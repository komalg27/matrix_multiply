* NGSPICE file created from multiply_komal.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlya_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_8 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlya_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

.subckt multiply_komal Clock Enable K[0] K[1] K[2] Result[0] Result[10] Result[11]
+ Result[12] Result[13] Result[14] Result[15] Result[16] Result[1] Result[2] Result[3]
+ Result[4] Result[5] Result[6] Result[7] Result[8] Result[9] X[0] X[1] X[2] X[3]
+ X[4] X[5] X[6] X[7] Z[0] Z[1] done reset vccd1 vssd1
XFILLER_67_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7957__A2 _2185_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5968__A1 _0998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7963_ _3103_ _3118_ _3132_ _3134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_54_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6914_ _2035_ _2036_ _2037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_51_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7894_ _2980_ _2987_ _3058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8657__CLK clknet_4_6_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7709__A2 _1701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6845_ _1779_ _1971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_52_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6776_ _1838_ _1903_ _1904_ _1905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_108_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8509__I1 _0112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8515_ _0084_ _3695_ _3711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5727_ _0823_ _0899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8134__A2 _1851_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6145__A1 _1146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8446_ _3633_ _3635_ _3640_ _3591_ _3638_ _3650_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5658_ _0827_ _0830_ _0831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_87_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7893__A1 _2974_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4609_ _3916_ _3931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8377_ _3546_ _3576_ _3577_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5589_ _0199_ _0345_ _0415_ _0386_ _0764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7328_ _2387_ _2450_ _2465_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6448__A2 _0063_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7645__A1 _0375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7259_ _2100_ _2390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6620__A2 _1755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5187__A2 _0354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4395__B1 _3478_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer7 _2189_ net40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_1
XFILLER_115_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7939__A2 _3106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4960_ _3809_ _4273_ _4274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4891_ _3840_ _4207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6630_ _1756_ _1765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__5178__A2 _3078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6561_ _1700_ _1701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4925__A2 _4239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8300_ _1094_ _1931_ _3496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5512_ _0686_ _0688_ _0689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6492_ _1569_ _1577_ _1636_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8231_ _3421_ _0103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5443_ _0611_ _0619_ _0620_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8162_ _3257_ _3344_ _3345_ _3346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5374_ _0494_ _0495_ _0551_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7113_ _2183_ _2231_ _2232_ _2234_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_99_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4325_ _2737_ _2745_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8093_ _3198_ _3235_ _3272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7044_ _1838_ _2164_ _2165_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5653__A3 _0414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8052__A1 _0564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8052__B2 _1734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7946_ _3113_ _3114_ _3115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4613__A1 _3813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7877_ _2974_ _2977_ _3041_ _3042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_58_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8355__A2 _0006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6828_ _1951_ _1953_ _1954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6759_ _1836_ _1853_ _1888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_17_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8107__A2 _1757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4403__I _3562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7866__A1 _0401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8429_ _3555_ _3561_ _3603_ _3632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_124_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7618__A1 _2742_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5234__I _0353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7094__A2 _2213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6841__A2 _1758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4852__A1 _3917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5580__A2 _0755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7857__A1 _0473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5144__I _0325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5090_ _0246_ _0272_ _0273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6832__A2 _1912_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7800_ _2933_ _2959_ _2960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_92_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5992_ _1150_ _1153_ _1154_ _1155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_64_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5399__A2 _0304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7731_ _2861_ _2866_ _2886_ _2887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_91_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4943_ _4256_ _4257_ _4258_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_91_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7662_ _0348_ _0352_ _2815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_32_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4874_ _4122_ _4190_ _4191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_18_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6613_ _1741_ _1749_ _1750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6899__A2 _1954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7593_ C\[0\]\[1\] _0184_ _2746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6544_ _1657_ _1659_ _1685_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6475_ _1451_ _1455_ _1620_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8214_ _3401_ _3403_ _3404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5426_ _0536_ _0543_ _0603_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8145_ _3274_ _3328_ _3329_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5357_ _3842_ _0413_ _0533_ _4169_ _0534_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7076__A2 _2128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8273__A1 _1672_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4308_ _2556_ _2567_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_8076_ _3251_ _3252_ _3253_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5288_ _0460_ _0466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7027_ _1529_ _1726_ _2148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4834__A1 A\[2\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4834__B2 _4077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4598__B1 _3196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7929_ _0577_ _1823_ _3096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6339__A1 _1477_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7000__A2 _2120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5562__A2 _4015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8687__D _0133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5314__A2 _4207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5865__A3 _4096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7067__A2 _2182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4825__A1 _4139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8016__A1 _3947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6290__A3 _0337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6578__A1 _0040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7619__I _1713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8319__A2 _2614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7790__A3 _2938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7782__C _3991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4590_ _3682_ _3909_ _3912_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6750__A1 _1824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8597__D _0042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6260_ _1306_ _1411_ _1330_ _1412_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5211_ _0391_ _0392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_83_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6191_ _1232_ _1236_ _1347_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5142_ _0309_ _0322_ _0323_ _0324_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8255__A1 _0607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5073_ _0228_ _0254_ _0255_ _0256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8007__A1 _3121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6569__A1 _3358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7230__A2 _1529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5975_ _1134_ _1137_ _1138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_80_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5241__A1 _3806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7714_ _0034_ _0925_ _1736_ _0002_ _2869_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4926_ _4238_ _4240_ _4241_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8694_ _0140_ clknet_4_7_0_Clock net30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5792__A2 _0891_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7645_ _0375_ _1758_ _2797_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4857_ _0043_ _4173_ _4174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7576_ _2721_ _2726_ _2730_ _2731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_4788_ _0056_ _4107_ _3907_ _4108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5544__A2 _0720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6527_ _1642_ _1669_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7297__A2 _2368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6458_ _1595_ _1602_ _1603_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5409_ _0524_ _0584_ _0586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6389_ _0337_ _1533_ _1535_ _1536_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7049__A2 _2147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8128_ _1371_ C\[0\]\[8\] _3228_ _3310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_62_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8059_ _3194_ _3198_ _3235_ _3236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_9_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7757__B1 _1702_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5783__A2 _0951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5535__A2 C\[2\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8485__A1 _0066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8485__B2 _0064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5299__A1 _4130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5299__B2 _0476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5471__A1 _0564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5223__A1 _0356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5760_ _0928_ _0929_ _0930_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8690__CLK clknet_4_5_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4711_ _4031_ _3863_ _4032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5691_ _0835_ _0836_ _0862_ _0863_ _0864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_7430_ _2511_ _2512_ _2575_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7515__A3 B\[1\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4642_ _3813_ _3964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5526__A2 _0654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7361_ _2282_ _2501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4573_ _3892_ _2836_ _3894_ _3895_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_128_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6312_ _1349_ _1353_ _1462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4501__I _3823_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7279__A2 _2013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7292_ _2424_ _2425_ _2426_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_115_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6243_ _1273_ _1395_ _1396_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8228__A1 _3351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6174_ _1307_ _1330_ _1331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_48_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8129__B _3310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5125_ _3271_ _0304_ _0306_ B\[2\]\[5\] _0307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__5332__I _0508_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5056_ _0193_ _0194_ _0239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_73_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5462__A1 _0422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8400__A1 _3462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7259__I _2100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5214__A1 _4275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5958_ _0675_ _0748_ _0821_ _1123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5765__A2 _0932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4909_ _4222_ _4223_ _4224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8677_ _0084_ clknet_4_12_0_Clock C\[3\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5889_ _0730_ _0742_ _1054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_107_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7628_ _2767_ _2780_ _2781_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_142_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6714__A1 _2492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7559_ _2712_ _2713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8563__CLK clknet_4_0_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5242__I _3831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5453__A1 _0564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6073__I _0607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5756__A2 _0049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6953__A1 _3562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4964__B1 _4216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6801__I _1927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5508__A2 _0609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6705__A1 _1247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4321__I _2695_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7130__A1 _0043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5152__I _0333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5444__A1 _0606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6930_ _4214_ _2053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6861_ _1981_ _1982_ _1986_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8600_ _0045_ clknet_4_9_0_Clock B\[1\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5812_ _4127_ _4144_ _0978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6792_ _1918_ _1919_ _1920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5743_ _0883_ _0884_ _0869_ _0915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_8531_ _0118_ _0073_ _3694_ _3725_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8536__I2 _0104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5674_ _0200_ _0467_ _0842_ _0847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
X_8462_ _3661_ _3790_ _0018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7413_ _2498_ _2555_ _2557_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4625_ _3946_ _3947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8393_ _0055_ _0015_ _3594_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7344_ _2422_ _2429_ _2482_ _2483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4556_ _3869_ _3878_ _3879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_102_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8586__CLK clknet_4_6_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7275_ _2335_ _2406_ _2407_ _2408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4487_ _3806_ _3809_ _3810_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6226_ _4173_ _0039_ _1380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7672__A2 _1716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5683__A1 _0854_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6157_ _1175_ _1186_ _1314_ _1315_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5108_ _0281_ _0290_ _0291_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6088_ _3842_ _0710_ _1248_ _1249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_44_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5435__A1 _4026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5435__B2 _0422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5039_ _0215_ _0221_ _0222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_2705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7188__A1 _2208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7360__A1 _2436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6163__A2 _3796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput20 net20 Result[13] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__7112__A1 _2184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput31 net31 Result[8] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__7663__A2 _1771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5674__A1 _0200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4477__A2 _3796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6218__A3 _0469_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5426__A1 _0536_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4316__I net15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8391__A3 _3500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4401__A2 _2755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6531__I _1672_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_118_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4410_ _3636_ _3646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5390_ _3978_ _0566_ _0567_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4341_ _2610_ _2362_ _2287_ _2908_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_67_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8458__I _0937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7103__A1 _2182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7060_ _3785_ _3866_ _1700_ _1998_ _2181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_98_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7654__A2 _2777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4468__A2 _3786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6011_ _1164_ _0337_ _1174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5417__A1 _0589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6706__I _3766_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7962_ _3121_ _3131_ _3132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6090__A1 _1249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6913_ _4227_ _2014_ _2036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7893_ _2974_ _3055_ _3057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6917__A1 _1973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6844_ _1960_ _1969_ _1970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_50_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6775_ _3971_ C\[1\]\[4\] _1904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7590__A1 _0033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7537__I _2689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8509__I2 _0082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8514_ _3707_ _3710_ _0139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5726_ _0206_ _0897_ _0898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8445_ _3623_ _3644_ _3648_ _3649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5657_ _0828_ _0829_ _0765_ _0830_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_108_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4608_ C\[3\]\[4\] _3826_ _3924_ _3929_ _3930_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5588_ _0760_ _0762_ _0763_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6696__A3 _1827_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8376_ _3549_ _3575_ _3576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_89_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7327_ _2464_ _0088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4539_ _3861_ _3862_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7272__I _2282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7645__A2 _1758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7258_ _2327_ _2340_ _2388_ _2389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5656__A1 _0386_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6209_ _1253_ _1256_ _1364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7189_ _2312_ _2314_ _2315_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_63_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_2_0_Clock_I clknet_3_1_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7948__A3 _3116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8601__CLK clknet_4_3_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6908__A1 _3776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7581__A1 _0920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4395__A1 _3391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4395__B2 B\[3\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7333__A1 _2400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer8 net42 net41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5895__A1 _0028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8133__I0 _3312_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5430__I _0408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6072__A1 _1057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4890_ _4197_ _4205_ _4206_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6375__A2 _1441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6560_ _3380_ _1698_ _1699_ A\[1\]\[0\] _3759_ _1700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_125_1171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5511_ _0027_ _0687_ _0688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6491_ _1575_ _1576_ _1635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5442_ _0614_ _0618_ _0619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8230_ _3343_ _3420_ _3421_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7875__A2 _3039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5886__A1 _0589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5373_ _0496_ _0550_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8161_ _3261_ _3330_ _3345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_47_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4324_ _2470_ _2737_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7112_ _2184_ _2186_ _2232_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8092_ _3262_ _3269_ _3270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7043_ _2163_ _2164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8624__CLK clknet_4_0_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5653__A4 _0823_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4861__A2 _4097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8052__A2 _0565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7945_ _3434_ _3110_ _1181_ _0566_ _1770_ _3114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4613__A2 _3934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7876_ _2989_ _3040_ _3041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_63_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6827_ _3499_ _1952_ _1953_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4377__A1 _3249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6758_ _1880_ _1886_ _1887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_6_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5709_ _0879_ _0880_ _0882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_109_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7315__A1 _2385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6689_ _1769_ _1773_ _1822_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8428_ _3607_ _3605_ _3609_ _3596_ _3631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7866__A2 _1252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8359_ _3462_ _0006_ _3558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7618__A2 _2743_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5629__A1 _0792_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5250__I _4159_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7306__A1 _2440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7857__A2 C\[0\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5868__A1 _1017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8647__CLK clknet_4_10_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6293__A1 _1433_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5991_ _0397_ _3867_ _1154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7793__A1 _0389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8471__I _3668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7730_ _2879_ _2885_ _2886_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_75_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4942_ _3912_ _4103_ _4257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7661_ _2809_ _2813_ _2814_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_127_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4873_ _4146_ _4149_ _4189_ _4190_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_21_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6612_ _3488_ _1748_ _1749_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7592_ _2742_ _2743_ _2744_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_119_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6543_ _1513_ _1514_ _1661_ _1684_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_119_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5571__A3 _0747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6474_ _1553_ _1618_ _1619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5859__A1 _3822_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8213_ _0633_ _2250_ _3403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5425_ _0536_ _0543_ _0602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_1250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8144_ _3296_ _3299_ _3327_ _3328_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5356_ _0353_ _0533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4307_ _2383_ _2556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_5287_ _0398_ _0461_ _0464_ _0465_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
X_8075_ _3153_ _3239_ _3252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6284__A1 _1184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5087__A2 _0243_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7026_ _2137_ _2145_ _2089_ _2146_ _2080_ _2147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_96_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4834__A2 _4078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8025__A2 _3128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7784__A1 _0435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4598__A1 _3919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7928_ _3992_ _0307_ _2237_ _3095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7859_ _3017_ _3018_ _3021_ _3022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_54_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5562__A3 _0537_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5314__A3 _0378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7067__A3 _2187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4825__A2 _4142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8016__A2 _0325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6578__A2 _1716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4589__A1 _3682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7790__A4 _2948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5305__A3 _0482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5210_ _0390_ _0391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__4513__A1 _3826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6190_ _1343_ _1345_ _1346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5141_ _0316_ _0321_ _0323_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_48_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8255__A2 _2123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5072_ _0231_ _0253_ _0255_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4816__A2 _4133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6569__A2 _3369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7766__A1 _2861_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7230__A3 _1975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5974_ _4131_ _1135_ _1136_ _0999_ _1137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_52_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5241__A2 _0415_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7713_ _0899_ _0001_ _0002_ _0925_ _2868_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4925_ C\[3\]\[3\] _4239_ _4240_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8693_ _0139_ clknet_4_5_0_Clock net29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7644_ _2766_ _2781_ _2795_ _2796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4856_ _4010_ _4173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7575_ _2701_ _2713_ _2728_ _2698_ _2729_ _2730_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_140_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4787_ _3899_ _4107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6526_ _1585_ _1642_ _1643_ _1668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_101_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6457_ _1601_ _1602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4504__A1 _3709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5408_ _0524_ _0584_ _0585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_88_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6388_ _1479_ C\[3\]\[13\] _1534_ _1535_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8127_ _3228_ _3227_ _3309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5339_ _0512_ _0472_ _0515_ _0516_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_47_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8058_ _3208_ _3219_ _3234_ _3235_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_87_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4807__A2 _4048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4409__I _3625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7009_ _2116_ _2129_ _2130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_99_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6009__A1 _4172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7757__A1 _0335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7757__B2 _0761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7509__A1 _2100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8182__A1 _3204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8485__A2 _3681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8237__A2 _3357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6248__A1 _1199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7996__A1 _3158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5471__A2 _0565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5223__A2 _0403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6420__A1 _1477_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4710_ _2878_ _4031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5690_ _0856_ _0860_ _0861_ _0863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7515__A4 _2665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4641_ _3961_ _3962_ _3796_ _3963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__6723__A2 _1832_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4572_ _3893_ _3894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7360_ _2436_ _2499_ _2500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_129_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6311_ _1458_ _1460_ _1461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7291_ _3968_ _2139_ _2425_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6487__A1 C\[2\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6242_ _1275_ _1272_ _1395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6173_ _1311_ _1329_ _1330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_97_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5124_ _0305_ _0306_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__7987__A1 _2760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5055_ _0149_ _0151_ _0164_ _0238_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_111_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5462__A2 _0393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8400__A2 _2665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5214__A2 _0374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5957_ _0675_ _0748_ _1122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4908_ _3801_ _3810_ _4223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8676_ _0083_ clknet_4_4_0_Clock C\[3\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5888_ _0693_ _0746_ _1052_ _1053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8164__A1 _3266_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4899__I _3757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7627_ _2768_ _2769_ _2779_ _2780_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_4839_ _4009_ _4157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__6714__A2 _1731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7911__A1 _3066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4725__A1 _3820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7558_ _2659_ _2711_ _2712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_107_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6509_ _1608_ _1610_ _1652_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7489_ _2542_ _2585_ _2638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4489__B1 _3391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5150__A1 _3982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5453__A2 _0565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6650__A1 _4157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6953__A2 _1848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8155__A1 _3052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4964__B2 _3774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7902__A1 _2994_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4716__A1 _3868_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7130__A2 _2250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_0_Clock_I Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6860_ _3931_ _1985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_1377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8394__A1 _3500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5811_ _4120_ _4191_ _0976_ _0977_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6791_ _3888_ _1865_ _1919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5747__A3 _0895_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8530_ _3724_ _0142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5742_ _0895_ _0912_ _0913_ _0914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8146__A1 _3270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8536__I3 _0089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8461_ _3661_ _0181_ _0017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5673_ _0802_ _0845_ _0846_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7412_ _2552_ _2553_ _2554_ _2555_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4624_ _2856_ _3946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_124_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8392_ _3590_ _3591_ _3571_ _3592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_102_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7343_ _2480_ _2428_ _2482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4555_ _3871_ _3874_ _3876_ _3877_ _3878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8449__A2 _1628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7274_ _2053_ _3873_ _1810_ _2404_ _2407_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_85_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4486_ _3808_ _3809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7121__A2 _2234_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6225_ _0716_ _0039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7672__A3 _2824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6156_ _1177_ _1312_ _1313_ _1314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_3_2_0_Clock_I clknet_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5107_ _0285_ _0286_ _0289_ _0290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6087_ _1247_ C\[2\]\[11\] _1248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_100_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6632__A1 _1760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5435__A2 _0364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5038_ _0024_ _0220_ _0221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input11_I X[6] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7188__A2 _2313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6935__A2 _2049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6989_ _2107_ _2108_ _2109_ _2110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_53_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8137__A1 _3301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8659_ _0128_ clknet_4_7_0_Clock C\[2\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7360__A2 _2499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6163__A3 _1319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5371__A1 _0528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput21 net21 Result[14] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_122_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput32 net32 Result[9] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__5123__A1 _2233_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8680__CLK clknet_4_7_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5674__A2 _0467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6871__A1 _2330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4477__A3 _3799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5426__A2 _0543_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5729__A3 _0825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8128__A1 _1371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4401__A3 _2764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4340_ _2589_ _2897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_126_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8300__A1 _1094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5163__I _0343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4468__A3 _3790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6010_ _0021_ _3998_ _1173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input3_I K[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6614__A1 _1738_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7961_ _3126_ _3130_ _3131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_54_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6090__A2 _1250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6912_ _2033_ _2034_ _2035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7892_ _2977_ _3041_ _3055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_74_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6843_ _1964_ _1968_ _1969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_63_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6917__A2 _2003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4928__A1 C\[3\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6774_ _1902_ _1903_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7590__A2 _1715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8513_ _0113_ _3708_ _3669_ _0128_ _3684_ _0083_ _3710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__8509__I3 _0127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5725_ _0896_ _0897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8444_ _3643_ _3647_ _3648_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5656_ _0386_ _0533_ _0829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5353__A1 _0397_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4607_ _3928_ _3929_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8375_ _3567_ _3574_ _3575_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5587_ _0206_ _0761_ _0762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7326_ _2456_ _2463_ _2464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_85_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4538_ _3260_ _2919_ _2298_ B\[3\]\[5\] _3861_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_105_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7257_ _2325_ _2342_ _2388_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4469_ _3775_ _3792_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_89_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5656__A2 _0533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6208_ _1361_ _1362_ _1363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6853__A1 _1895_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7188_ _2208_ _2313_ _2229_ _2226_ _2314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_86_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6139_ _1006_ _1296_ _1297_ _1153_ _1298_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6605__A1 _3746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4417__I _3701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8358__A1 _1673_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_6_0_Clock_I clknet_3_3_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6908__A2 _3004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7030__A1 _3894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8052__C _3960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7581__A2 _1772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4395__A2 _2405_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5592__A1 _0489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer9 _3604_ net42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5344__A1 _0492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6687__A4 _1793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5895__A2 _0445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6844__A1 _1960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8576__CLK clknet_4_1_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7021__A1 _2138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5583__A1 _0021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5158__I _0022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5510_ _0444_ _0687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6490_ _1481_ _1572_ _1633_ _1634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8521__A1 _3715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5441_ _0615_ _0616_ _0617_ _0618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_86_1421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8160_ _3261_ _3330_ _3344_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5372_ _0494_ _0495_ _0549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7111_ _2184_ _2186_ _2231_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7088__A1 _0059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4323_ _2460_ _2717_ _2727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_113_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8091_ _3266_ _3268_ _3269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_141_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6835__A1 _3864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7042_ _2075_ _2076_ _3100_ _2163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8037__B1 _3112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4310__A2 net8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5621__I _0476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7260__A1 _1768_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7944_ _0651_ _1714_ _3112_ _3113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_82_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7260__B2 _2313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7875_ _2992_ _3039_ _3040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__7012__A1 _2072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6452__I _1528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6826_ _1930_ _1952_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6757_ _1884_ _1885_ _1886_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_91_1171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5708_ _0879_ _0880_ _0881_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_104_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6688_ _1774_ _1797_ _1820_ _1821_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5326__A1 _3315_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8427_ _3589_ _3628_ _3629_ _3630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5639_ _0452_ _0585_ _0813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_128_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8358_ _1673_ _3556_ _3557_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7309_ _2430_ _2444_ _2445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8289_ _3427_ _3484_ _3485_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_120_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6627__I _1762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4852__A3 _4169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8599__CLK clknet_4_3_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7003__A1 _3229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4368__A2 net6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8503__A1 _3692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7306__A2 _2441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5317__A1 _3315_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5868__A2 _1033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6817__A1 _3889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6293__A2 _1443_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5990_ _3862_ _3293_ _1153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7793__A2 _1894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4941_ _4234_ _4254_ _4255_ _4256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7660_ _2811_ _2812_ _2813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4872_ _4165_ _4188_ _4189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6611_ _1747_ _1748_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5556__A1 _3615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7591_ _0436_ _1826_ _2743_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6542_ _1664_ _1682_ _1683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_53_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6473_ _1555_ _1552_ _1618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6221__B _1375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8212_ _3398_ _3399_ _3400_ _3401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5859__A2 _3824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5424_ _0546_ _0583_ _0600_ _0601_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8143_ _3320_ _3325_ _3327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_86_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5355_ _0440_ _0530_ _0531_ _0532_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_82_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4306_ _2492_ _2513_ _2534_ A\[3\]\[3\] _2545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_8074_ _3155_ _3250_ _3251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5286_ _3983_ C\[2\]\[4\] _0464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_87_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7025_ _2085_ _2088_ _2146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6284__A2 _4080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6036__A2 _0178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7233__A1 _0514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7784__A2 _2257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7927_ _3091_ _3093_ _3094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_71_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7858_ _3019_ _1770_ _3020_ _1181_ _3021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_58_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6809_ _1874_ _1923_ _1935_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7789_ _2946_ _1771_ _1972_ _2947_ _2948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_71_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5562__A4 _0533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8497__B1 _3695_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5314__A4 _0036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8016__A3 _1755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7224__A1 _3969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7775__A2 _2932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5786__A1 _0919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6092__I _1252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7916__I _3005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8614__CLK clknet_4_3_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8488__B1 _3669_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4340__I _2589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5710__A1 _0870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5140_ _0316_ _0321_ _0322_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_123_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6266__A2 _1300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7463__A1 _2550_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6267__I _1295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5071_ _0231_ _0253_ _0254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_29_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8482__I _3675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6569__A3 _1707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5777__A1 _0024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5973_ _0982_ _1000_ _1136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7230__A4 _2087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7712_ _2860_ _2865_ _2866_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4924_ _3928_ _4239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8692_ _0138_ clknet_4_5_0_Clock net28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7643_ _2767_ _2780_ _2795_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5529__A1 _0703_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4855_ _4172_ _0043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8191__A2 _2045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6730__I _1699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7574_ _2694_ _2714_ _2729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4786_ _3902_ _3906_ _4106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_105_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6525_ _1666_ _1667_ _0078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6456_ _1596_ _1599_ _1600_ _1601_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5407_ _0546_ _0583_ _0584_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5701__A1 _0847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4504__A2 _3766_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6387_ _0795_ _1534_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8126_ _3303_ _3307_ _3308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5338_ _0514_ C\[2\]\[6\] _0515_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_115_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8057_ _3224_ _3233_ _3234_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5269_ _0442_ _0446_ _0447_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_60_1210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7008_ _2118_ _2128_ _2129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_75_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4807__A3 _4064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6009__A2 _4062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4283__A4 _2287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7757__A2 _0752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5768__A1 _0016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4425__I _3747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8637__CLK clknet_4_0_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5256__I _0434_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5940__A1 _4072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6248__A2 _1202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7996__A2 _3160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6956__B1 _1990_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6971__A3 _2093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8173__A2 _3357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4640_ _3936_ _3962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_129_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7920__A2 _3035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6723__A3 _1854_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4571_ _3358_ net12 _3893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4734__A2 _4048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6310_ _1342_ _1458_ _1459_ _1460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_128_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7290_ _3816_ _2281_ _2424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6241_ _1121_ _1124_ _1393_ _1394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6487__A2 _1630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6172_ _1315_ _1328_ _1329_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_135_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5123_ _2233_ _2254_ _3747_ _2287_ _0305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_84_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7987__A2 _2103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5054_ _0192_ _0235_ _0236_ _0237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5998__A1 _1017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5214__A3 _0377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5956_ _0866_ _0964_ _0967_ _0749_ _1121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_90_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4907_ _4217_ _4219_ _4221_ _4222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8675_ _0082_ clknet_4_5_0_Clock C\[3\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5887_ _0695_ _0745_ _1052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_51_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8164__A2 _3268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7626_ _2770_ _2777_ _2778_ _2779_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_4838_ _4154_ _4082_ _4155_ _4156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7911__A2 _3075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7557_ _2709_ _2710_ _2711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4725__A2 _4045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5922__A1 _4218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4769_ _3542_ _4089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5922__B2 _3773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6508_ _1592_ _1593_ _1651_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7488_ _2544_ _2584_ _2637_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7675__A1 _2819_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6439_ _1583_ _1584_ _1585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4489__A1 A\[2\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5150__A2 _3892_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8109_ _3088_ _3287_ _3288_ _3190_ _3289_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7978__A2 _0962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6650__A2 _1783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4413__A1 _0056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4964__A2 _4220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7466__I _2501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6166__A1 _1184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7363__B1 _2152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6705__A3 _1723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5913__A1 _4026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8538__S0 _3678_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7666__A1 _0823_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7130__A3 _2141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8091__A1 _3266_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5810_ _4122_ _4190_ _0976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6790_ _1916_ _1917_ _1918_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4404__A1 _2794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5741_ _0910_ _0911_ _0913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8460_ _0937_ _3981_ _0046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5672_ _0843_ _0844_ _0794_ _0845_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7411_ _1372_ C\[1\]\[12\] _2552_ _2554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_15_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4623_ C\[3\]\[5\] _3929_ _3939_ _3945_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4707__A2 _3849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8391_ _0055_ _0015_ _3500_ _3591_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_135_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7342_ _2359_ _2480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4554_ _3864_ _3877_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7657__A1 _0752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7273_ _3873_ _1810_ _2404_ _2053_ _2406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4485_ _3807_ _3808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6224_ _1037_ _0037_ _1379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_131_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7409__A1 _3999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6155_ _1180_ _1182_ _1185_ _1313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5106_ _0288_ _0289_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6086_ _0456_ _1247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8156__B _3331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5037_ _3903_ _0220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_3_6_0_Clock_I clknet_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8385__A2 _3541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6396__A1 _1526_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6988_ _2025_ _2094_ _2109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6935__A3 _2057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4946__A2 _4260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5939_ _1102_ _1103_ _1104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6148__A1 _1167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8658_ _0127_ clknet_4_6_0_Clock C\[2\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6699__A2 _1793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7609_ _2759_ _2760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_120_1421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8589_ _0034_ clknet_4_2_0_Clock B\[0\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput22 net22 Result[15] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_107_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6871__A2 _1707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8128__A2 C\[0\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6139__A1 _1006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6139__B2 _1153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_114_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8300__A2 _1931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7960_ _3127_ _3128_ _3129_ _3130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_82_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6911_ _3903_ _1952_ _2034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7891_ _3053_ _3041_ _3054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8367__A2 _3566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6842_ _1965_ _1966_ _1967_ _1968_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_74_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6773_ _1846_ _1849_ _2674_ _1902_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4928__A2 _4242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8512_ _3686_ _3708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5724_ _0343_ _0896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5655_ _3875_ _0364_ _0828_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8443_ _3626_ _3622_ _3647_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4606_ _3927_ _3928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8374_ _3568_ _3573_ _3574_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5353__A2 _0529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5586_ _0317_ _0761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_4_13_0_Clock_I clknet_3_6_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7325_ _2457_ _2462_ _2463_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4537_ _3859_ _3860_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7256_ _2316_ _2376_ _2386_ _2387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4468_ _3778_ _3786_ _3790_ _3791_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_132_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_1411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6207_ _1259_ _1265_ _1362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7187_ _3026_ _1929_ _2313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4399_ _2470_ _3531_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_58_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4864__A1 _3948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8055__A1 _3230_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6138_ _1150_ _1154_ _1297_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7502__C _2602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6605__A2 _3748_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6069_ _1090_ _1091_ _1231_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_3227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4616__A1 _3822_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5041__A1 _0180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4433__I _3755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5592__A2 _0199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7869__A1 _0924_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6541__A1 _1590_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5344__A2 _0497_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8294__A1 _3452_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8046__A1 _0487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5280__A1 _0457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6823__I _1864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7021__A2 _2140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5032__A1 _0026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5583__A2 _0757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8521__A2 _3716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5440_ _4061_ _0423_ _0617_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6532__A1 _3434_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4543__B1 _3562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5371_ _0528_ _0547_ _0520_ _0519_ _0502_ _0548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_103_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5174__I _0354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7110_ _2226_ _2229_ _2230_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4322_ _2706_ _2717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7088__A2 _2120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8090_ _3092_ _3267_ _3183_ _3180_ _3268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_99_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7041_ _1018_ _1840_ _2161_ _2162_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__6835__A2 _1882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4846__A1 _4156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8037__A1 _0716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8037__B2 _3976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4518__I _3840_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7260__A2 _2390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7943_ _3423_ _3110_ _3112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6733__I _1863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7874_ _3008_ _3012_ _3038_ _3039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_63_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6825_ _1948_ _1950_ _1951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_50_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6771__A1 _3832_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6756_ _3786_ _1791_ _1885_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8670__CLK clknet_4_4_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5707_ _0841_ _0846_ _0880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_109_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6687_ _1719_ _1819_ _1794_ _1793_ _1820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__7564__I _2718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8600__D _0045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8426_ _3610_ _3612_ _3629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_104_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5638_ _0789_ _0810_ _0811_ _0812_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5326__A2 _0461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7866__A4 _1736_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5569_ _0695_ _0745_ _0746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8357_ _1528_ C\[0\]\[13\] _3556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8276__A1 _0718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7308_ _2433_ _2443_ _2444_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8288_ _3428_ _3483_ _3484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7239_ _2364_ _2368_ _2369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_77_106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8028__A1 _0384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5262__A1 _2695_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7003__A2 _2123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5259__I _0315_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6514__A1 _1595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5317__A2 _0493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6817__A2 _0012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4828__A1 _4124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5253__A1 _3413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4940_ _4252_ _4253_ _4255_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8693__CLK clknet_4_5_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4871_ _4167_ _4187_ _4188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_2890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6610_ _1746_ _1747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7590_ _0033_ _1715_ _2742_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5556__A2 _0529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6541_ _1590_ _1616_ _1650_ _1682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6472_ _1590_ _1616_ _1617_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6505__A1 _1619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5423_ _0548_ _0582_ _0600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_118_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8211_ _0630_ _2275_ _3400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5859__A3 _4179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5354_ _0310_ _0408_ _0531_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8142_ _3323_ _3324_ _3325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4305_ _2524_ _2534_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_82_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8073_ _3238_ _3250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5285_ _0374_ _0458_ _0462_ _0463_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7024_ _2074_ _2078_ _2145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6284__A3 _4176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5492__A1 _0625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6036__A3 _0300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5244__A1 _0422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7926_ _3069_ _3092_ _3093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5795__A2 _0962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7857_ _0473_ C\[0\]\[6\] _3020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6808_ _1871_ _1932_ _1933_ _1934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5547__A2 _0709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7788_ _0387_ _0388_ _2947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_23_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6739_ _1866_ _1867_ _1868_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5807__I _4107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8497__A1 _0087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8497__B2 _0117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8409_ _3564_ _3566_ _3611_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4507__B1 _3829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8566__CLK clknet_4_0_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5483__A1 C\[2\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6027__A3 _1189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7224__A2 _0003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5786__A2 _0932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8185__B1 _2102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8488__A1 _0068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8488__B2 _0070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5070_ _0210_ _0234_ _0252_ _0253_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_111_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5226__A1 _3848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5972_ _0060_ _0030_ _1135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5777__A2 _0048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7711_ _2862_ _2863_ _2864_ _2865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_4923_ _3997_ _3818_ _4238_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8691_ _0137_ clknet_4_5_0_Clock net27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7642_ _2783_ _2782_ _2793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6726__A1 _1760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4854_ _3948_ _3936_ _4172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5529__A2 _0704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4785_ _3912_ _4103_ _4104_ _4105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7573_ _2694_ _2714_ _2728_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_119_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6524_ _1647_ _1648_ _1665_ _1667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8589__CLK clknet_4_2_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6455_ _1598_ C\[3\]\[14\] _1596_ _1600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5406_ _0548_ _0582_ _0583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_47_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6386_ _1531_ _1533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5701__A2 _0873_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4504__A3 _3804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8125_ _3305_ _3306_ _3307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5337_ _0513_ _0514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_130_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5362__I _0353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5268_ _0201_ _0445_ _0446_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8056_ _3225_ _3232_ _3233_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_130_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7007_ _2125_ _2127_ _2128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_112_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5199_ _0349_ _0380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_116_1492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7757__A3 _2911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5768__A2 _0925_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6965__A1 _4157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7909_ _2760_ _2203_ _3074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6717__A1 _2599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7238__B _2367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4441__I _3753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7142__A1 _2252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7996__A3 _3166_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5208__A1 _0387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6956__A1 _4003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6956__B2 _4088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8532__B _3708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4351__I _3004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4570_ _3067_ _3892_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6240_ _1120_ _1272_ _1273_ _1393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_115_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5695__A1 _0020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6171_ _1318_ _1327_ _1328_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5182__I _0362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5122_ _0303_ _0304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__7436__A2 _2581_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5053_ _0196_ _0197_ _0236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5998__A2 _1033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4526__I _2963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5214__A4 _0384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5955_ _1116_ _1119_ _1120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4422__A2 net8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4906_ _3791_ _4220_ _4221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8674_ _0081_ clknet_4_4_0_Clock C\[3\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5886_ _0589_ _0593_ _0692_ _0691_ _0684_ _1051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_16_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7625_ C\[0\]\[2\] _0184_ _2778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4837_ _4046_ _4068_ _4155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6175__A2 _1331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7372__A1 _1538_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7556_ _2702_ _2703_ _2708_ _2710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
Xclkbuf_4_14_0_Clock clknet_3_7_0_Clock clknet_4_14_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4768_ _4087_ _4088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4725__A3 _3937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5922__A2 _0647_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6507_ _1649_ _1615_ _1650_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7124__A1 _2147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4699_ _3944_ _4019_ _4020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7487_ _2596_ _2635_ _2636_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_135_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6438_ _1558_ _1560_ _1582_ _1584_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__7675__A2 _2823_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5686__A1 _0854_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6369_ _1515_ _1516_ _1517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5150__A3 _0331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7427__A2 _2487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8108_ _3186_ _3189_ _3288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_103_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5438__A1 _3615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8039_ _3211_ _3212_ _3213_ _3214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8604__CLK clknet_4_1_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6938__A1 _1989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5610__A1 _0780_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4413__A2 _0030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7363__A1 _1319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5267__I _0444_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6166__A2 _4079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7363__B2 _1164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6705__A4 _1781_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4716__A3 _4036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5913__A2 _0409_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8538__S1 _3719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7666__A2 _1783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5730__I _0901_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8091__A2 _3268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6929__A1 _4133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4404__A2 _2836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6561__I _1700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5740_ _0910_ _0911_ _0912_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5671_ _0342_ _0498_ _0793_ _0795_ _0844_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__7354__A1 _2367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7410_ C\[1\]\[12\] _3929_ _2553_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4622_ _3914_ _3942_ _3943_ _3944_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8390_ _3569_ _3570_ _3590_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4553_ _3875_ _3876_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7341_ _2477_ _2478_ _2479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7106__A1 _4112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7657__A2 _1702_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4484_ B\[1\]\[0\] _3754_ _3380_ _3756_ _3701_ _3807_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_7272_ _2282_ _2404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5668__A1 _0776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6223_ _1377_ _1378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8627__CLK clknet_4_8_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7409__A2 _2404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6154_ _1180_ _1182_ _1185_ _1312_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_140_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6736__I _1740_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5105_ _0246_ _0272_ _0287_ _0288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6085_ _0374_ _1099_ _1101_ _1246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4684__C _3938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6093__A1 _0541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5036_ _3882_ _0024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5840__A1 _0800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6987_ _2025_ _2094_ _2108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_53_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8603__D _0048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5938_ _0800_ _0710_ _1101_ _3976_ _1103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_80_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8657_ _0126_ clknet_4_6_0_Clock C\[2\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7345__A1 _3877_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5869_ _4069_ _0020_ _4068_ _1035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_107_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7608_ _0467_ _2759_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8588_ _0033_ clknet_4_2_0_Clock B\[0\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7539_ _2682_ _2688_ _2690_ _2691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5815__I _3315_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7648__A2 _1748_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput23 net23 Result[16] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_135_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6320__A2 _1358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5123__A3 _3747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5831__A1 _4156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6381__I _4085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8128__A3 _3228_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7336__A1 _2411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5725__I _0896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6847__B1 _1910_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4873__A2 _4149_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8064__A2 _3137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7811__A2 _2961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5822__A1 _0973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6910_ _1966_ _2030_ _2032_ _2033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7890_ _2977_ _3053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6841_ _4200_ _1758_ _1967_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6772_ _1896_ _1900_ _1901_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_143_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8511_ _0098_ _3681_ _3707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5723_ _4073_ _0032_ _0895_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8442_ _3645_ _0108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7878__A2 _3042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5654_ _0824_ _0825_ _0826_ _0827_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5889__A1 _0730_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4605_ _3423_ _3926_ _3927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8373_ _3569_ _3570_ _3571_ _3573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_5585_ _3876_ _0315_ _0760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7324_ _2458_ _2459_ _2461_ _2462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_89_1272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4536_ _3858_ _3859_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7255_ _2320_ _2375_ _2386_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_131_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4467_ _3789_ _3790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6206_ _1245_ _1258_ _1361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6853__A3 _1908_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7186_ _2310_ _2311_ _2312_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4398_ _3510_ _0056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4864__A2 _3824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6137_ _0419_ _1295_ _1296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7802__A2 _2961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6068_ _1090_ _1091_ _1230_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5813__A1 _4124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4616__A2 _3936_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5019_ _0203_ _4227_ _0204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4714__I _4034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5592__A3 _0345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7869__A2 _2257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8046__A2 _2250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5280__A2 C\[2\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4624__I _2856_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7021__A3 _2141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5032__A2 _0207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7309__A1 _2430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6780__A2 _1908_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6532__A2 _1671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5370_ _0492_ _0497_ _0547_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4543__B2 _2919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4321_ _2695_ _2706_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8285__A2 _3452_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7670__I _0403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7040_ _3925_ _2159_ _2161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4846__A2 _4163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8037__A2 _2771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7942_ C\[0\]\[7\] _3110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7873_ _3010_ _3025_ _3036_ _3038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_51_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7012__A3 _2090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6824_ _3218_ _1949_ _1950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6220__A1 _1374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6755_ _1878_ _1881_ _1883_ _1884_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_56_1282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6771__A2 _1899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5706_ _0872_ _0875_ _0876_ _0878_ _0879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_104_1214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6686_ _1795_ _1819_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8425_ _3610_ _3612_ _3628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_104_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5637_ _0808_ _0809_ _0811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5326__A3 _0474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4534__A1 _3413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8356_ _3521_ _3523_ _3554_ _3555_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5568_ _0698_ _0724_ _0744_ _0745_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_88_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7307_ _2439_ _2442_ _2443_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_132_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4519_ _3841_ _3842_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8276__A2 _1987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8287_ _3430_ _3482_ _3483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5499_ _0598_ _0676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6287__A1 _4066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7238_ _2365_ _2366_ _2367_ _2368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_137_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4837__A2 _4068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8028__A2 _1252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7169_ _2291_ _2293_ _2294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_98_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7787__A1 _0379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5262__A2 _0319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4444__I _3766_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8200__A2 _3325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8519__C _3714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5253__A2 _3467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4870_ _4175_ _4186_ _4187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_2891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6540_ _1619_ _1621_ _1665_ _1617_ _1681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_119_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6471_ _1612_ _1615_ _1616_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_101_1409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6505__A2 _1621_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8210_ _1181_ _3398_ _3399_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5422_ _0588_ _0598_ _0599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5859__A4 _4180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8141_ _0899_ _2614_ _3128_ _3324_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_99_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5353_ _0397_ _0529_ _0530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4304_ _2254_ _2276_ _2524_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8072_ _3248_ _0130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5284_ _0461_ _0462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7023_ _2136_ _2143_ _2144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_101_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6284__A4 _1322_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7769__A1 _0308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7233__A3 _2156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5244__A2 _0423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7925_ _0314_ _1862_ _3092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6992__A2 _2093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7856_ _0504_ _0505_ _3019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6807_ _1872_ _1924_ _1933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7787_ _0379_ _0381_ _2946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5547__A3 _0723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4999_ _0184_ _0185_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8611__D _0056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6738_ _1818_ _1856_ _1867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_143_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8497__A2 _3693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6669_ _1803_ _0087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8408_ _3596_ _3609_ _3610_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4507__B2 _3770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8339_ _3428_ _3483_ _3537_ _3538_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5180__A1 _4072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4439__I _3761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5483__A2 _3860_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6680__A1 _0202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6680__B2 _3510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4443__B1 _3196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4994__A1 _3979_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8185__A1 _0750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8185__B2 _0051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5219__B _3946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8488__A2 _3687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7999__A1 _3121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8660__CLK clknet_4_14_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6564__I _1703_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5971_ _0980_ _0060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4434__B1 _2341_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7710_ _0335_ _0896_ _2237_ _2864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4922_ _4222_ _4223_ _4237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8690_ _0136_ clknet_4_5_0_Clock net26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7641_ _2784_ _2782_ _2792_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4853_ _4068_ _4170_ _4171_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_60_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7923__A1 _2926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4812__I _3293_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4737__A1 _3955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7572_ _2722_ _2725_ _2726_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_119_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4784_ _4022_ _4102_ _4104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_18_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6523_ _1647_ _1648_ _1665_ _1666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_118_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6454_ _1598_ C\[3\]\[14\] _1534_ _1599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_31_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5405_ _0559_ _0563_ _0581_ _0582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__5162__A1 _2816_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5162__B2 B\[2\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6385_ _1528_ C\[3\]\[13\] A\[2\]\[6\] _0047_ _1532_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_8124_ _0487_ _1986_ _3306_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5336_ _3854_ _0513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8055_ _3230_ _3231_ _3232_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_88_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5267_ _0444_ _0445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6662__A1 _1793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7006_ _3888_ _2126_ _2127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5198_ _3853_ _2578_ _0346_ B\[0\]\[4\] _0379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_99_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_10_0_Clock clknet_3_5_0_Clock clknet_4_10_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__8606__D _0051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6965__A2 _2087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7908_ _3071_ _3072_ _3073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8167__A1 _3274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7839_ _2998_ _2999_ _3000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_54_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7914__A1 _3012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6717__A2 _1848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8683__CLK clknet_4_12_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6653__A1 _3402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5208__A2 _0388_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6956__A2 _1770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7905__A1 _2928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4719__A1 _4025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5695__A2 _0757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6170_ _1321_ _1325_ _1326_ _1327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_124_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5121_ _3727_ _2276_ _2556_ _0303_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_111_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5052_ _0196_ _0197_ _0235_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6947__A2 _1993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4958__A1 _4270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5954_ _0678_ _1117_ _1118_ _1119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4905_ _3794_ _4002_ _3799_ _4220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_8673_ _0080_ clknet_4_4_0_Clock C\[3\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5885_ _1050_ _0086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8556__CLK clknet_4_2_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7624_ _2772_ _2774_ _2776_ _2777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_4836_ _4044_ _4074_ _4154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_107_1459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7372__A2 _0005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7555_ _2702_ _2703_ _2708_ _2709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4767_ _3925_ _4087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6506_ _1612_ _1649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7486_ _2598_ _2634_ _2635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4698_ _3988_ _4018_ _4019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8321__A1 _3518_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5135__A1 _3819_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6437_ _1558_ _1560_ _1582_ _1583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_115_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6368_ _0062_ _3900_ _3646_ _0063_ _1516_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_103_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8107_ _0577_ _1757_ _3287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5319_ _4072_ _0393_ _0496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6299_ _1409_ _1449_ _1450_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5438__A2 _0363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8038_ _0718_ _1736_ _3213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4646__B1 _3967_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6938__A2 _2001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7060__A1 _3785_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4949__A1 _0027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5610__A2 _0782_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4452__I _2856_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6166__A3 _4176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7363__A2 _1999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8312__A1 _3461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5283__I _0460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4401__B A\[3\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5429__A2 _0558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4637__B1 _3954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8379__A1 _3495_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8379__B2 _3493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8579__CLK clknet_4_6_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6929__A2 _1882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4404__A3 _3572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4362__I _3122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5670_ _0199_ _0498_ _0842_ _0843_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8551__A1 _3704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7354__A2 _2437_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5365__A1 _0541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4621_ _3930_ _3941_ _3943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7340_ _2409_ _2413_ _2478_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4552_ _3122_ _3875_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8303__A1 _0445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7271_ _2401_ _2402_ _2403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4483_ _3805_ _3806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6865__A1 _3982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6222_ _1366_ _1376_ _1377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_48_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6153_ _1172_ _1308_ _1310_ _1311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5104_ _0270_ _0271_ _0287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6084_ _1243_ _1108_ _1244_ _1245_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7290__A1 _3816_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6093__A2 _0037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5035_ _0188_ _0190_ _0219_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_85_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5840__A2 _3873_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6986_ _2022_ _2107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7593__A2 _0184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5937_ _0800_ _0710_ _1101_ _1102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_53_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8656_ _0125_ clknet_4_6_0_Clock C\[2\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5868_ _1017_ _1033_ _1034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8542__A1 _3693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7345__A2 _2123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7607_ _0945_ _0010_ _2757_ _2758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4819_ _4135_ _4137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8587_ _0032_ clknet_4_1_0_Clock B\[0\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5799_ _0965_ _0967_ _0968_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7538_ _2650_ _2681_ _2690_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5108__A1 _0281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7469_ _2613_ _2615_ _2617_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_134_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5659__A2 _0830_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6856__A1 _2492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput24 net24 Result[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_89_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5123__A4 _2287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6608__A1 _3792_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4447__I _3749_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5292__B1 _0464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5831__A2 _4163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5595__A1 _3772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5278__I _4089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8533__A1 _0088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7336__A2 _2473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6847__A1 _3962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6847__B2 _1893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6075__A2 _1235_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6840_ _2460_ _1811_ _1966_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6771_ _3832_ _1899_ _1900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4306__B A\[3\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8510_ _3706_ _0138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5722_ _0894_ _0032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5338__A1 _0514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8441_ _3624_ _3644_ _3645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5653_ _4275_ _3871_ _0414_ _0823_ _0826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4604_ _3925_ _3926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8372_ _3446_ _3569_ _3501_ _3498_ _3571_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_5584_ _0754_ _0758_ _0759_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_129_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7323_ _2301_ _2378_ _2461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4535_ _3760_ _3856_ _3857_ _3858_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_117_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6838__A1 _1961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7254_ _2382_ _2384_ _2385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4466_ A\[2\]\[2\] _3787_ _2826_ _3788_ _3789_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_132_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6205_ _1359_ _1360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7185_ _2223_ _2243_ _2311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4397_ _3499_ _3510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6136_ _4137_ _1295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4864__A3 _4179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6067_ _1089_ _1229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5018_ _2889_ _0203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4616__A3 _3937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8614__D _0059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5577__A1 _0207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6969_ _2064_ _2091_ _2092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8515__A1 _0084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5592__A4 _0415_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8639_ _0095_ clknet_4_2_0_Clock C\[1\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5501__A1 _0588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7006__A1 _3888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5032__A3 _4117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8617__CLK clknet_4_9_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4640__I _3936_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6532__A3 _1673_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4543__A2 _2930_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4320_ _2685_ _2695_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_114_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7493__A1 _2536_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input1_I Enable vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7245__A1 _2320_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7941_ _3107_ _3108_ _3109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_110_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4815__I _3867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7872_ _3028_ _3031_ _3035_ _3036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_51_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5559__A1 _0574_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6823_ _1864_ _1949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6220__A2 C\[2\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6754_ _4202_ _1882_ _1883_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5705_ _0848_ _0877_ _0878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__7347__B _2485_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6251__B _1335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6685_ _1813_ _1817_ _1818_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4550__I _3872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5636_ _0808_ _0809_ _0810_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8424_ _3500_ _3594_ _3592_ _3627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_12_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8355_ _3518_ _0006_ _3524_ _3554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5567_ _0727_ _0743_ _0744_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4534__A2 _2794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7306_ _2440_ _2441_ _2442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4518_ _3840_ _3841_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8286_ _3435_ _3481_ _3482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5498_ _0451_ _0673_ _0674_ _0675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7237_ _1178_ C\[1\]\[9\] _2155_ _2139_ _2367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__7484__A1 _2611_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6287__A2 _0755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8609__D _0054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4449_ _3771_ _3772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7168_ _2111_ _2193_ _2292_ _2293_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_113_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8028__A3 _3104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7236__A1 _4090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6119_ _1278_ _0119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7099_ _2216_ _2217_ _2218_ _2219_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_59_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7787__A2 _0381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5291__I _0468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4635__I _3934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5253__A3 _0380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8551__B _3686_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6850__I _1975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6470_ _1509_ _1549_ _1614_ _1615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7702__A2 _2778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5421_ _0594_ _0597_ _0598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4516__A2 _2982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8140_ _3321_ _3322_ _3323_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5352_ _0314_ _0529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4303_ _2503_ _2513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8071_ _0965_ _0967_ _3248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_141_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5283_ _0460_ _0461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7022_ _2137_ _2142_ _2143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_87_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7769__A2 _1701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7233__A4 _1903_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7924_ _0363_ _1929_ _3091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7855_ _0514_ C\[0\]\[6\] _0569_ net43 _3018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_51_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6806_ _1872_ _1924_ _1932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7786_ _2937_ _2944_ _2945_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4998_ _4242_ _0184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6737_ _0057_ _0008_ _1749_ _1759_ _1866_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_17_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4280__I net2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6668_ _1800_ _1802_ _1803_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5619_ _3973_ C\[2\]\[2\] _0793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8407_ _3605_ _3608_ _3609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4507__A2 _3769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6599_ _1735_ _1736_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8338_ _3430_ _3482_ _3537_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5180__A2 _0360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7457__A1 _2179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8269_ _3462_ _0003_ _3399_ _3463_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_65_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7209__A1 _2053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5483__A3 _3928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6680__A2 _0010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4455__I _3777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4443__B2 _3765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4994__A2 _0179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8185__A2 _2013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6196__A1 _0054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5943__A1 _1105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7696__A1 _0903_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6845__I _1779_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7620__A1 _0539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5970_ _1132_ _1133_ _1134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4434__B2 _3756_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4921_ _4235_ _4236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_92_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7640_ _2791_ _0117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4852_ _3917_ _3762_ _4169_ _4170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7923__A2 _3088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7571_ _2707_ _2723_ _2724_ _2725_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4783_ _4022_ _4102_ _4103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4737__A2 _4007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5196__I _0376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6522_ _1650_ _1664_ _1665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8501__S _3668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6453_ _1597_ _1598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5404_ _0516_ _0573_ _0580_ _0581_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_118_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6384_ _1531_ _0047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8123_ _0509_ _1899_ _3305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7439__A1 _2544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5335_ net37 _0512_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_86_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8054_ _0633_ _3104_ _3231_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5266_ _0443_ _0444_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7005_ _2102_ _2126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5197_ _0377_ _0378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5622__B1 _0466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7907_ _0903_ _2579_ _3072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4976__A2 _0153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8622__D _0110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7838_ _2236_ _0307_ _2911_ _2999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_54_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7914__A2 _3038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5925__A1 _0541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4728__A2 _3963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7769_ _0308_ _1701_ _2926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_32_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6653__A2 _1707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4664__A1 _3970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4967__A2 _4204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6169__A1 _3961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7905__A2 _3069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5120_ _0302_ _0085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8094__A1 _3198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5051_ _0217_ _0232_ _0233_ _0234_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6575__I _1713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4655__A1 _3973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5953_ _0681_ _0747_ _1118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4958__A2 _4271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4904_ _4218_ _3809_ _4219_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5884_ _1047_ _1049_ _1050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8672_ _0072_ clknet_4_4_0_Clock C\[3\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7623_ _0333_ net34 _2776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4835_ _4150_ _4151_ _4152_ _4057_ _4058_ _4153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_60_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6580__A1 _1479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7554_ _2666_ _2704_ _2707_ _2708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4766_ _3983_ C\[3\]\[7\] _3964_ _4085_ _4086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_140_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6505_ _1619_ _1621_ _1617_ _1648_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7485_ _2607_ _2633_ _2634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4697_ _3996_ _4006_ _4017_ _4018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__8321__A2 _0005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6436_ _1561_ _1581_ _1582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6367_ _1419_ _0063_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8085__A1 _3184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8106_ _3283_ _3285_ _3286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5318_ _3773_ _0401_ _0495_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6298_ _1410_ _1448_ _1449_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8617__D _0062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5249_ _0373_ _0427_ _0428_ _0429_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8037_ _0716_ _2771_ _3112_ _3976_ _3212_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_103_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4646__B2 _3765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4949__A2 _3240_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_8_0_Clock clknet_3_4_0_Clock clknet_4_8_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_12_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7899__A1 _2983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6166__A4 _1322_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5374__A2 _0495_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8650__CLK clknet_4_11_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4885__A1 _3056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6395__I _1541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4637__A1 _3825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4637__B2 _3958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7051__A2 _2057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4643__I _3964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8551__A2 _0123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4620_ _3930_ _3941_ _3942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5365__A2 _0423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4551_ _3873_ _3874_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5474__I _0648_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8303__A2 _2579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7270_ _3864_ _1928_ _2402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4482_ _3804_ _3805_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6221_ _1370_ _1373_ _1375_ _1376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8067__A1 _3052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6152_ _4173_ _0045_ _1174_ _1310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5103_ _0161_ _0170_ _0286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_112_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7814__A1 _2909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6083_ _1100_ _1102_ _1103_ _1244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5034_ _0191_ _0198_ _0217_ _0218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7290__A2 _2281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6985_ _2016_ _2104_ _2105_ _2106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4553__I _3875_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5936_ _3983_ C\[2\]\[10\] _1101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4800__A1 _4107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8673__CLK clknet_4_4_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8655_ _0117_ clknet_4_12_0_Clock C\[2\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5867_ _1024_ _1032_ _1033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7606_ _0375_ _1748_ _2757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4818_ _3111_ _4135_ _4136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8586_ _0031_ clknet_4_6_0_Clock A\[3\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5798_ _0966_ _0820_ _0967_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_124_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7537_ _2689_ _0092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4749_ _3955_ _4070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7468_ _2613_ _2615_ _2616_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_107_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput25 net25 Result[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_135_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6856__A2 _1731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6419_ _1488_ _1565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7399_ _2479_ _2489_ _2541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4619__A1 _3939_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5292__A1 _4207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5292__B2 _0469_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8230__A1 _3343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4463__I _3785_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5595__A2 _0354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8533__A2 _3681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4555__B1 _3876_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5294__I _0460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8297__A1 _3441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6847__A2 _1972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4638__I _3946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8696__CLK clknet_4_13_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5469__I _0568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_0 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6770_ _1897_ _1898_ _1899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5721_ _0336_ _0334_ _0894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8440_ _3626_ _3643_ _3644_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5338__A2 C\[2\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5652_ _0489_ _0033_ _0825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4603_ net15 _3925_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5583_ _0021_ _0757_ _0758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8371_ _0687_ _2103_ _3570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7322_ _2301_ _2378_ _2459_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4534_ _3413_ _2794_ _3369_ _2836_ _3857_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_50_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6838__A2 _1963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7253_ _2309_ _2315_ _2384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4465_ _3779_ _3445_ _2513_ _3788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_85_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4849__A1 _3970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6204_ _1357_ _1358_ _1359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7184_ _2225_ _2242_ _2310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4396_ _3488_ _3499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6135_ _1292_ _1293_ _1294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4548__I _3870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4864__A4 _4180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6066_ _1070_ _1080_ _1228_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8460__A1 _0937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5274__A1 _0340_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5017_ _3904_ _0202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5577__A2 _0752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6968_ _2068_ _2073_ _2090_ _2091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_53_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5919_ _0709_ _0723_ _1084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6899_ _1945_ _1954_ _2021_ _2022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8515__A2 _3695_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8630__D _0104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5329__A2 _0505_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8638_ _0087_ clknet_4_9_0_Clock C\[1\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8569_ _0014_ clknet_4_3_0_Clock A\[1\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8279__A1 _0037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8569__CLK clknet_4_3_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6829__A2 _1954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4458__I _3780_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6673__I _1765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8203__A1 _3311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7006__A2 _2126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5289__I _0466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_5_0_Clock clknet_0_Clock clknet_3_5_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_41_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7190__A1 _2309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5752__I _0359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6583__I _1721_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7940_ _0392_ _2250_ _3108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7871_ _3032_ _3033_ _3034_ _3035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__5008__A1 _4270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6822_ _1881_ _1946_ _1947_ _1948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5559__A2 _0537_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6756__A1 _3786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6220__A3 B\[2\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6753_ _1739_ _1882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5704_ _0871_ _0873_ _0843_ _0877_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6684_ _1815_ _1816_ _1817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8423_ _3613_ _3616_ _3626_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5635_ _0486_ _0521_ _0454_ _0809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_117_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8354_ _3550_ _3552_ _3553_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5566_ _0730_ _0742_ _0743_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_30_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4534__A3 _3369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7305_ _4085_ _1962_ _2441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4517_ _3838_ _3839_ _3775_ _3840_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_105_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5497_ _0587_ _0672_ _0674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8285_ _3438_ _3452_ _3480_ _3481_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_132_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7236_ _4090_ C\[1\]\[9\] _3974_ _2366_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6287__A3 _4179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4448_ _3768_ _3769_ _2341_ _3770_ _3771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_104_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4278__I net3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4379_ _3304_ _3315_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7167_ _2114_ _2192_ _2292_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_99_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8028__A4 _1907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6118_ _1274_ _1277_ _1278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7098_ _2135_ _2170_ _2218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5247__A1 _0406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8625__D _0113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6049_ _1069_ _1113_ _1211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_41_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6747__A1 _1832_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4758__B1 _4078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4741__I _4061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7475__A2 _0185_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5486__A1 _3133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8424__A1 _3500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8551__C _3741_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4651__I _3972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5420_ _0595_ _0596_ _0597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5713__A2 _0884_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5351_ _0492_ _0497_ _0528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_57_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4302_ _2383_ _2503_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_8070_ _3247_ _0115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5282_ _0430_ _0304_ _0306_ _0459_ _0460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_114_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5477__A1 _4071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7021_ _2138_ _2140_ _2141_ _2142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_59_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6674__B1 _1743_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5229__A1 _3133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7923_ _2926_ _3088_ _3090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_97_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7854_ _3013_ _3014_ _3016_ _3017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_23_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6805_ _1931_ _0013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7785_ _2938_ _2942_ _2943_ _2944_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__5401__A1 _4033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4997_ _4270_ _0180_ _0182_ _0183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4561__I _3883_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6736_ _1740_ _0008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5952__A2 _0747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7154__A1 _0513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6667_ _1722_ _1751_ _1801_ _1802_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8406_ _3606_ _3607_ _3608_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5618_ _0465_ _0470_ _0792_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5704__A2 _0873_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6598_ _1732_ _1734_ _1735_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8337_ _3489_ _3535_ _3536_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5549_ _0725_ _0618_ _0726_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5392__I _0568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7457__A2 _2390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8268_ _0632_ _3462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7219_ _2260_ _2261_ _2347_ _2348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8199_ _3301_ _3319_ _3387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8607__CLK clknet_4_1_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7209__A2 _2282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5483__A4 _0658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4443__A2 _3764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4471__I _3793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7932__A3 _3098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5943__A2 _1106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6499__A3 _1641_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7696__A2 _1811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6120__A2 _1192_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6959__A1 _3950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7620__A2 _2771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4434__A2 _3754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4920_ _4224_ _4225_ _4235_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_3391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6082__B _1100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4851_ _4168_ _4169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7570_ _1673_ _2707_ _2723_ _2724_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4782_ _4041_ _4101_ _4102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4737__A3 _3831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6521_ _1651_ _1653_ _1663_ _1664_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__7136__A1 _3817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6452_ _1528_ _1597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5403_ _0575_ _0578_ _0579_ _0580_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_6383_ _4070_ _1530_ _1531_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8122_ _0392_ _3302_ _3303_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4370__A1 _3196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5334_ _0507_ _0510_ _0511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_47_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8053_ _3227_ _3226_ _3228_ _3230_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5265_ _0325_ _0443_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7004_ _2122_ _2124_ _2125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_9_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5196_ _0376_ _0377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7611__A2 _0008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5622__B2 _2717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7906_ _3001_ _3068_ _3070_ _3071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7837_ _0326_ _1823_ _2998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_19_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4291__I net4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7768_ _2870_ _2877_ _2925_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5925__A2 _0488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6719_ _1847_ _1850_ _1851_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7699_ _2850_ _2851_ _2852_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_138_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_4_0_Clock clknet_3_2_0_Clock clknet_4_4_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_59_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5861__A1 _0513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6681__I _1808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7118__A1 _4214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5050_ _0191_ _0198_ _0233_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_69_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4655__A2 _3976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5604__A1 _3814_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5952_ _0681_ _0747_ _1117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_18_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4903_ _4071_ _4218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8671_ _0065_ clknet_4_4_0_Clock C\[3\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5883_ _4261_ _0301_ _1048_ _1049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7357__A1 _1247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7622_ _2773_ _1980_ _2774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4834_ A\[2\]\[7\] _4078_ _3894_ _4077_ _4152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__5000__I _0185_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7553_ _2666_ _2705_ _2707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_14_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4765_ _4084_ _3764_ _4060_ _3765_ _4085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__6580__A2 C\[1\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6504_ _1590_ _1616_ _1647_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7484_ _2611_ _2632_ _2633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4696_ _4008_ _4011_ _4016_ _4017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_105_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6435_ _1563_ _1580_ _1581_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_106_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6366_ _1513_ _1514_ _1515_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_1_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8105_ _3267_ _3284_ _3285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5317_ _3315_ _0493_ _0494_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6297_ _1413_ _1447_ _1448_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6096__A1 _1254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8036_ _0716_ _1715_ _3112_ _3211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5248_ _0406_ _0426_ _0428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4646__A2 _3764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5179_ _0358_ _0359_ _3990_ _0360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_96_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7596__A1 _0375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8633__D _0107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7060__A3 _1700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4885__A2 _3089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6676__I _1808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6087__A1 _1247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7823__A2 _2981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5834__A1 _3849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4924__I _3928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7339__A1 _2403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6011__A1 _1164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5755__I _0903_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4573__A1 _3892_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4550_ _3872_ _3873_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4481_ _3802_ _3750_ _3744_ _3803_ _3804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__7511__A1 _2659_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6220_ _1374_ C\[2\]\[12\] B\[2\]\[7\] _0981_ _1375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_83_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5704__B _0843_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6151_ _1309_ _0045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5102_ _0282_ _0283_ _0284_ _0285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6082_ _1102_ _1103_ _1100_ _1243_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5825__A1 _4149_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5033_ _0210_ _0213_ _0216_ _0217_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7578__A1 _0048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5589__B1 _0415_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6984_ _2019_ _2095_ _2105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5935_ _0342_ _1099_ _0712_ _1100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_80_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4800__A2 _4117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8654_ _0071_ clknet_4_4_0_Clock C\[2\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5866_ _1026_ _1030_ _1031_ _1032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__6002__A1 _1164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7605_ _2756_ _0071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4817_ _4034_ _4135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8585_ _0030_ clknet_4_6_0_Clock A\[3\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5797_ _0814_ _0819_ _0966_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5665__I _0377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4564__A1 _3837_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7536_ _2682_ _2688_ _2689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4748_ _3917_ _4069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7467_ _1538_ _2614_ _2615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7502__A1 _2603_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4679_ _3997_ _3825_ _3999_ _4000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6418_ _1490_ _1492_ _1564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput26 net26 Result[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_7398_ _2483_ _2488_ _2540_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4867__A2 _4183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8628__D _0116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6349_ _1464_ _1498_ _1499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5816__A1 _0980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8019_ _3188_ _3191_ _3192_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_29_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5292__A2 _0467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7569__A1 _1688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6241__A1 _1121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4555__A1 _3871_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4555__B2 _3877_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8297__A2 _3451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8541__I0 _0121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4858__A2 _4174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_3_1_0_Clock clknet_0_Clock clknet_3_1_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_95_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5720_ _0892_ _0893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_62_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5651_ _3871_ _0050_ _0823_ _4275_ _0824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4546__A1 _3865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4602_ _3918_ _3923_ _3924_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8370_ _0055_ _0014_ _3569_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5582_ _0436_ _0757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_129_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7321_ _2291_ _2293_ _2458_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4533_ _3854_ _3467_ _2764_ _3855_ _3856_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_102_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7252_ _2312_ _2314_ _2382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4464_ _3402_ _2352_ _3748_ _3782_ _3787_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_131_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6203_ _1262_ _1263_ _1230_ _1358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_89_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7183_ _0220_ _0015_ _2211_ _2309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4395_ _3391_ _2405_ _3478_ B\[3\]\[0\] _3488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_98_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6134_ _1149_ _1156_ _1293_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6065_ _1083_ _1112_ _1226_ _1227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8460__A2 _3981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5016_ _0201_ _0025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8640__CLK clknet_4_0_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8480__B _3679_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6967_ _2074_ _2078_ _2089_ _2090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_5918_ _1073_ _1082_ _1083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_107_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6898_ _1944_ _2020_ _2021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8637_ _0067_ clknet_4_0_0_Clock C\[1\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5849_ _4181_ _4183_ _4185_ _1015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7723__A1 _2870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8568_ _0013_ clknet_4_3_0_Clock A\[1\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7519_ _2664_ _2669_ _2670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_120_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8279__A2 _3302_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8499_ _0102_ _3666_ _3697_ _0072_ _3698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_68_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7115__I _1753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4474__I _3078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7962__A1 _3121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7718__C _2236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7714__A1 _0034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4649__I _3854_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8663__CLK clknet_4_14_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4384__I net5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7870_ _0435_ _2562_ _3034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5008__A2 _0180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6821_ _0980_ _1761_ _1824_ _1947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_93_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7953__A1 _3013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6756__A2 _1791_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6752_ _2449_ _1765_ _1881_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6220__A4 _0981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5429__B _0605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5703_ _0200_ _0838_ _0876_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6683_ _0211_ _1748_ _1763_ _1812_ _1816_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__7705__A1 _2819_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8422_ _3622_ _3623_ _3624_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5634_ _0790_ _0806_ _0807_ _0808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7181__A2 _2288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8353_ _0481_ _0007_ _3527_ _3552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5565_ _0735_ _0741_ _0742_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_121_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4534__A4 _2836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7304_ _3917_ _2350_ _2440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4516_ _3067_ _2982_ _2631_ _3839_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_89_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8284_ _3455_ _3479_ _3480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5496_ _0587_ _0672_ _0673_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8130__A1 _0514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4559__I _3870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7235_ _3957_ _2139_ _2365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4447_ _3749_ _3770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6287__A4 _1437_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6692__A1 _1768_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7166_ _2198_ _2290_ _2291_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_63_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4378_ _3293_ _3304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6117_ _1275_ _1276_ _1277_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6774__I _1902_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7097_ _2190_ _2217_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6048_ _1209_ _1210_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8197__A1 _3368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7999_ _3121_ _3131_ _3170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__7944__A1 _0651_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6747__A2 _1854_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8641__D _0097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4758__A1 _3819_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4758__B2 A\[2\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8686__CLK clknet_4_13_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4469__I _3775_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6683__A1 _0211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4997__A1 _4270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8188__A1 _3992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7163__A2 _2248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5350_ _0412_ _0525_ _0526_ _0527_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8112__A1 _3287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4379__I _3304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4301_ _2481_ _2492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5281_ B\[2\]\[0\] _0459_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_64_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7020_ _3980_ _1971_ _2141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6674__A1 _2897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5477__A2 _0571_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6674__B2 A\[1\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6594__I _1709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5229__A2 _0409_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4328__B A\[3\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7922_ _3960_ _0325_ _2050_ _3088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_64_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7853_ _0387_ _0388_ _1847_ _1850_ _1753_ _3016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_82_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8559__CLK clknet_4_8_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7926__A1 _3069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6804_ _1930_ _1931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7784_ _0435_ _2257_ _2943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4996_ _3979_ _3799_ _4150_ _0181_ _0182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5401__A2 _0577_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6735_ _1865_ _0012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6666_ _1738_ _1750_ _1801_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5617_ _0776_ _0779_ _0791_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8405_ _3553_ _3563_ _3607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6597_ _3078_ _1733_ _1734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_30_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8336_ _3492_ _3534_ _3535_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5548_ _0614_ _0725_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8103__A1 _0343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4289__I net2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8267_ _3459_ _3460_ _3461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5479_ _0576_ _0656_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7218_ _2258_ _2259_ _2347_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8198_ _3366_ _3385_ _3386_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_59_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8636__D _0066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7149_ _2270_ _2271_ _2272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4428__B1 _3745_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4979__A1 _4222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output26_I net26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7917__A1 _3000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4752__I _4072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_4_0_0_Clock clknet_3_0_0_Clock clknet_4_0_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_1478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8342__A1 _3424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6679__I _1811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5156__A1 _0336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7853__B1 _1847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4927__I _3927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6959__A2 _1971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8701__CLK clknet_4_13_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4850_ _3804_ _4168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5395__A1 _3953_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4781_ _4043_ _4100_ _4101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6520_ _1655_ _1662_ _1663_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_18_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7136__A2 _2257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8333__A1 _3512_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5147__A1 _0324_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6451_ _4152_ _1533_ _1596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5698__A2 _3870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5402_ C\[2\]\[7\] _4242_ _0579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6382_ _1529_ _1530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8121_ _2077_ _3302_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5333_ _3921_ _0509_ _0510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4370__A2 _2405_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6647__A1 _0457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8052_ _0564_ _0565_ _1732_ _1734_ _3960_ _3228_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_5264_ _0410_ _0439_ _0441_ _0442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_115_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4658__B1 _3572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7003_ _3229_ _2123_ _2124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5195_ _0375_ _0376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_68_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5870__A2 _4174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7905_ _2928_ _3069_ _3070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4572__I _3893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7836_ _2938_ _2995_ _2996_ _2944_ _2937_ _2997_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_34_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5386__A1 _0511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7767_ _2866_ _2922_ _2923_ _2924_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4979_ _4222_ _4223_ _4245_ _0165_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_6718_ _1849_ _1850_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8324__A1 _1672_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7698_ _2759_ _1865_ _2851_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6649_ _3972_ C\[1\]\[2\] _3975_ _1784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_69_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8319_ _0481_ _2614_ _3517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6638__A1 _3786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5861__A2 C\[3\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7063__A1 _3821_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5613__A2 _0786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4482__I _3804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7366__A2 _2506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6169__A3 _4096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5377__A1 _3604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7118__A2 _2164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6877__A1 _1979_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6629__A1 _0211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5301__A1 _3531_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4657__I _3978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4655__A3 C\[3\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7054__A1 _3991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5604__A2 _0383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5951_ _1051_ _1115_ _1116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_111_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4902_ _3774_ _4216_ _4217_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_55_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8670_ _0064_ clknet_4_4_0_Clock C\[3\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5882_ _4194_ _4260_ _1048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7357__A2 C\[1\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5368__A1 _0528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7621_ _0922_ _0923_ _2773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4833_ _4057_ _4058_ _4151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_107_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5907__A3 _0740_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7552_ C\[1\]\[15\] _1630_ _2705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4764_ B\[1\]\[7\] _4084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8306__A1 _3497_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6503_ _1646_ _0123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6580__A3 _0040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7483_ _2620_ _2630_ _2632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4695_ _4012_ _4015_ _4016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6868__A1 _3957_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6434_ _1564_ _1579_ _1580_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_140_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6365_ _3900_ _1419_ _1514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5540__A1 _4273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8104_ _0314_ _2011_ _3284_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5316_ _0376_ _0493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6296_ _1425_ _1446_ _1447_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_27_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5172__B _3593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8035_ _3113_ _3114_ _3116_ _3210_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4567__I _3888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6096__A2 _1255_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5247_ _0406_ _0426_ _0427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5178_ _3456_ _3078_ _0350_ _0359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7045__A1 _2160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7596__A2 _1704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7060__A4 _1998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8545__A1 _3719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7819_ _2914_ _2915_ _2978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6859__A1 _4001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5531__A1 _0661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7284__A1 _2358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6087__A2 C\[2\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5834__A2 _3615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7036__A1 _1372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7587__A2 _0951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7339__A2 _2408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6011__A2 _0337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5770__A1 _0937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4573__A2 _2836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4480_ A\[2\]\[4\] _3803_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5522__A1 _0637_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6150_ _4158_ _4003_ _1309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5101_ _0267_ _0269_ _0284_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4387__I _2233_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6081_ _1240_ _1241_ _1242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_48_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5032_ _0026_ _0207_ _4117_ _0215_ _0216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_111_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7027__A1 _1529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7578__A2 _0008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5589__A1 _0199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6983_ _2019_ _2095_ _2104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5589__B2 _0386_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5934_ _0657_ _1099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8527__A1 _0131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8527__B2 _0086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8653_ _0070_ clknet_4_4_0_Clock C\[2\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5865_ _4045_ _4067_ _4096_ _1031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__4850__I _3804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7604_ _0944_ _0952_ _2756_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4816_ _3859_ _4133_ _4134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5796_ _0866_ _0964_ _0965_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8584_ _0029_ clknet_4_4_0_Clock A\[3\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7750__A2 _2887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5761__A1 _0928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7535_ _2646_ _2684_ _2687_ _2688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4747_ _4066_ _4067_ _3950_ _4068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_135_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7466_ _2501_ _2614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4678_ _3998_ _3999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7502__A2 _2604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6417_ _1472_ _1496_ _1562_ _1563_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6777__I _1905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7397_ _2537_ _2538_ _2539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput16 net16 Result[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput27 net27 Result[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_1_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6348_ _1468_ _1497_ _1498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_116_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4297__I _2438_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6279_ _1323_ _1324_ _1326_ _1430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_103_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5816__A2 _0981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8018_ _3186_ _3189_ _3190_ _3191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_69_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8644__D _0100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6241__A2 _1124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4555__A2 _3874_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8541__I1 _0076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7257__A1 _2325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7009__A1 _2116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5991__A1 _0397_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8592__CLK clknet_4_10_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4670__I _3991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5650_ _0822_ _0823_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7732__A2 _2887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4601_ _3762_ _3922_ _3817_ _3923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4546__A2 _3868_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5581_ _0756_ _0021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7320_ _2295_ _2294_ _2296_ _2379_ _2457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_2
X_4532_ A\[3\]\[0\] _3855_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7251_ _2381_ _0101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4463_ _3785_ _3786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6202_ _1233_ _1357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7182_ _2215_ _2305_ _2306_ _2307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4394_ _3434_ _2352_ _3445_ _3467_ _3478_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_28_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6133_ _1152_ _1155_ _1292_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7799__A2 _2958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6064_ _1086_ _1111_ _1226_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5015_ _0200_ _0201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6471__A2 _1615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7221__I _2164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6966_ _2080_ _2085_ _2088_ _2089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_81_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5917_ _1077_ _1081_ _1082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6897_ _1955_ _2020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8636_ _0066_ clknet_4_1_0_Clock C\[1\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5848_ _4181_ _4183_ _4185_ _1014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_107_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7723__A2 _2877_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5734__A1 _3882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8567_ _0012_ clknet_4_0_0_Clock A\[1\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5779_ C\[2\]\[0\] _0947_ _0948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7518_ _2666_ _2668_ _2669_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8498_ _3679_ _3678_ _3697_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8639__D _0095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7449_ _2576_ _2581_ _2595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7239__A1 _2364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4755__I _3818_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7411__A1 _1372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5973__A1 _0982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5586__I _0317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4490__I _3812_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7714__A2 _0925_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4528__A2 _3850_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6150__A1 _4158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8522__S0 _3683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4464__A1 _3402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6820_ _4202_ _1740_ _1761_ _4195_ _1946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_63_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7953__A2 _3014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6751_ _1769_ _1878_ _1879_ _1827_ _1880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_50_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5702_ _0848_ _0874_ _0875_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6682_ _4116_ _0009_ _1763_ _1814_ _1815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_52_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7705__A2 _2823_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8421_ _3581_ _3618_ _3619_ _3623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_104_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5716__A1 _0835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5633_ _0804_ _0805_ _0807_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5564_ _0736_ _0737_ _0740_ _0741_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_8352_ _2665_ _0007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7303_ _2367_ _2437_ _2439_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4515_ _3037_ _3048_ _2534_ A\[3\]\[4\] _3838_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_8283_ _3458_ _3461_ _3477_ _3479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_144_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5495_ _0599_ _0671_ _0672_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_89_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6141__A1 _3874_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7234_ _2279_ _2283_ _2363_ _2364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4446_ _3735_ _3769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_104_216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7165_ _2201_ _2289_ _2290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__6692__A2 _1747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4377_ _3249_ _3282_ _3100_ _3293_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6116_ _1120_ _1125_ _1276_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7096_ _2135_ _2170_ _2216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4575__I _3896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6047_ _1207_ _1208_ _1209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8197__A2 _3384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7998_ _3168_ _3109_ _3117_ _3169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_1627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4758__A2 _4077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6949_ _2069_ _2070_ _2071_ _2072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8619_ _0068_ clknet_4_1_0_Clock C\[0\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8510__I _3706_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4930__A2 _4244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5486__A3 _0662_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7880__A1 _2839_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6683__A2 _1748_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4997__A2 _0180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7796__I _2955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8188__A2 _0576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7148__B1 _0004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7163__A3 _2286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8630__CLK clknet_4_10_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4300_ _2470_ _2481_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5280_ _0457_ C\[2\]\[3\] _0458_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_86_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6674__A2 _1742_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7623__A1 _0333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7921_ _3084_ _3085_ _3086_ _3087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_110_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7852_ _0379_ _0381_ _2871_ _2872_ _3100_ _3014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_93_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7926__A2 _3092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6803_ _1929_ _1930_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5937__A1 _0800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7783_ _2939_ _2940_ _2942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4995_ _4002_ _0181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6734_ _1864_ _1865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6665_ _1799_ _1800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7154__A3 _2652_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8404_ _3555_ _3561_ _3606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5616_ _0773_ _0783_ _0790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6596_ _1707_ _1733_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_121_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8335_ _3493_ _3533_ _3534_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_117_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5547_ _0707_ _0709_ _0723_ _0724_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_118_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8103__A2 _2099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8266_ _3405_ _3410_ _3460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5478_ _0653_ _0654_ _0655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7862__A1 _3023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7217_ _2264_ _2344_ _2345_ _2346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4429_ B\[1\]\[2\] _3752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_120_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8197_ _3368_ _3384_ _3385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7148_ _1530_ _1826_ _0004_ _4069_ _2271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7079_ _2132_ _2191_ _2199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4428__A1 _3718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6968__A3 _2090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8652__D _0094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8653__CLK clknet_4_4_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5156__A2 _0337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7853__A1 _0387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7853__B2 _1850_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4667__A1 _3758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6644__B _3760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8562__D _0007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8030__A1 _0822_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5919__A1 _0709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4780_ _4050_ _4065_ _4099_ _4100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_61_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6592__A1 _4157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5395__A2 _0571_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6450_ _1537_ _1539_ _1532_ _1595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5401_ _4033_ _0577_ _0578_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5698__A3 _4239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6895__A2 _2006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6381_ _4085_ _1529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_103_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5332_ _0508_ _0509_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8120_ _3224_ _3233_ _3300_ _3301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5263_ _0316_ _0440_ _0441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7844__A1 _3000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8051_ _3926_ _3226_ _3227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4658__A1 B\[1\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4658__B2 _3783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7002_ _2013_ _2123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5194_ _3797_ _0311_ _0312_ B\[2\]\[1\] _0375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_5_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5014__I _0199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7904_ _3792_ _0317_ _3002_ _3069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_52_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8676__CLK clknet_4_4_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8021__A1 _3177_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7835_ _2942_ _2943_ _2996_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7766_ _2861_ _2886_ _2923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_71_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4978_ _4238_ _4240_ _0164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6717_ _2599_ _1848_ _1849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4594__B1 _3802_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7697_ _2849_ _2811_ _2850_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_71_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6648_ net38 _1783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__6335__A1 _4161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5689__A3 _0861_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6579_ _1688_ C\[1\]\[0\] _1630_ _1718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8088__A1 _3179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8318_ _3514_ _3515_ _3516_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8088__B2 _3177_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8647__D _0089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6638__A2 _1772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8249_ _3439_ _3440_ _3441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5377__A2 _0376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8315__A2 _3475_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6877__A2 _1989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4888__A1 _4201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8079__A1 _3158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8557__D _0002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6629__A2 _0009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5301__A2 _2786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8699__CLK clknet_4_13_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7054__A2 _2993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8251__A1 _0053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5950_ _1053_ _1114_ _1115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_53_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4901_ _4070_ _4213_ _4215_ _4216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_80_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5881_ _0972_ _1046_ _1047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_61_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7357__A3 _0476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7620_ _0539_ _2771_ _2772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4832_ _3807_ _4150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__6565__A1 _0208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7551_ C\[1\]\[15\] _0947_ _2704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4763_ _4075_ _4082_ _4083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6502_ _1644_ _1645_ _1646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6580__A4 _1715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7482_ _2623_ _2629_ _2630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4694_ _4014_ _4015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6868__A2 _1725_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6433_ _1568_ _1578_ _1579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_88_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6364_ _1421_ _1513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5540__A2 _0716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8103_ _0343_ _2099_ _3283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5315_ _0490_ _0404_ _0491_ _0492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6295_ _1428_ _1445_ _1446_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8034_ _3107_ _3108_ _3209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5246_ _0412_ _0418_ _0425_ _0426_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_29_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4500__B1 _3797_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5177_ _3853_ _2578_ _0346_ B\[0\]\[1\] _0358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_68_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5056__A1 _0193_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4583__I _3636_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8545__A2 _0092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7818_ _2921_ _2975_ _2976_ _2977_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_51_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7749_ _2847_ _2902_ _2903_ _2904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6859__A2 _4150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8481__A1 _3660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8233__A1 _3343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7036__A2 C\[1\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5770__A2 _0181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4573__A3 _3894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5522__A2 _0638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5100_ _0267_ _0269_ _0283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6080_ _1093_ _1110_ _1241_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5286__A1 _3983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5031_ _0214_ _0208_ _0215_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7027__A2 _1726_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5038__A1 _0024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6786__A1 _0202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6982_ _2103_ _0015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5589__A2 _0345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6250__A3 _1335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5933_ _1096_ _0722_ _1097_ _1098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_81_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8652_ _0094_ clknet_4_11_0_Clock C\[1\]\[16\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5864_ _1028_ _1029_ _1030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7603_ _2754_ _0065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4815_ _3867_ _4133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6002__A3 _1019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8583_ _0028_ clknet_4_4_0_Clock A\[3\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5795_ _0893_ _0962_ _0963_ _0964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7534_ _2686_ _2687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4746_ _3795_ _4067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4564__A3 _3879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7465_ _1419_ _2579_ _2613_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4677_ _3934_ _3998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6416_ _1493_ _1495_ _1562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_rebuffer10_I _1713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6710__A1 _0513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7396_ _2474_ _2519_ _2538_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput17 net17 Result[10] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput28 net28 Result[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__4578__I _3899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6347_ _1472_ _1496_ _1497_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_66_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6278_ _1316_ _1317_ _1429_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_102_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5277__A1 _0396_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8017_ _2236_ _0308_ _3002_ _3190_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_102_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5229_ _3133_ _0409_ _0410_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_88_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5202__I _0382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8660__D _0129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5201__A1 _0379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7129__I _1899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5872__I _1037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6701__A1 _1374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5268__A1 _0201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8206__A1 _0632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6768__A1 _3542_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5440__A1 _4061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8570__D _0015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5991__A2 _3867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4600_ _3921_ _3922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5743__A2 _0884_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6940__A1 _1974_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5580_ _3822_ _0755_ _0756_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4531_ _3853_ _3854_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_117_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7250_ _2379_ _2380_ _2381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_89_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4462_ B\[1\]\[2\] _3781_ _2826_ _3784_ _3785_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_102_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6201_ _1239_ _1267_ _1355_ _1356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4398__I _3510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7181_ _2219_ _2288_ _2306_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4393_ _3456_ _3467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6132_ _1160_ _1289_ _1290_ _1291_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6063_ _1061_ _1224_ _1225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5014_ _0199_ _0200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6759__A1 _1836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6965_ _4157_ _2087_ _2088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5431__A1 _2717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5916_ _1070_ _1080_ _1081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_81_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6896_ _1939_ _2017_ _2018_ _2019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8635_ _0109_ clknet_4_11_0_Clock C\[0\]\[16\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5847_ _4165_ _4188_ _1012_ _1013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7184__A1 _2225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8566_ _0011_ clknet_4_0_0_Clock A\[1\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5734__A2 _0903_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5778_ _0186_ _0947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7517_ _1533_ _2152_ _2667_ _2668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4729_ _4048_ _4049_ _3986_ _4050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8497_ _0087_ _3693_ _3695_ _0117_ _3696_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_120_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7448_ _2594_ _0090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5498__A1 _0451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7379_ _2474_ _2519_ _2520_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7239__A2 _2368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8655__D _0117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6998__A1 _2031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5670__A1 _0199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5422__A1 _0588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7714__A3 _1736_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5489__A1 _0661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6150__A2 _4003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8565__D _0010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8522__S1 _3704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4464__A2 _2352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7938__B1 _1903_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5413__A1 _0398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4681__I _3823_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6750_ _1824_ _1825_ _1879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5701_ _0847_ _0873_ _0874_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6681_ _1808_ _1814_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_108_1377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8420_ _3588_ _3617_ _3622_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5632_ _0804_ _0805_ _0806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6913__A1 _4227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8351_ _3520_ _3526_ _3550_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5563_ _0738_ _0617_ _0739_ _0740_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7302_ _2434_ _2435_ _2436_ _2437_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4514_ _3811_ _3835_ _3836_ _3837_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8282_ _3473_ _3476_ _3477_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5494_ _0601_ _0670_ _0671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7233_ _0514_ C\[1\]\[8\] _2156_ _1903_ _2363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__8529__S _3714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4445_ A\[2\]\[2\] _3768_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6141__A2 _0981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5017__I _3904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7164_ _2215_ _2219_ _2288_ _2289_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_119_1462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4376_ _3067_ _3271_ _2631_ _3282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_99_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6115_ _1116_ _1119_ _1275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4856__I _4010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7095_ _2205_ _2214_ _2215_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_112_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6046_ _0689_ _1064_ _1208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5652__A1 _0489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7997_ _3022_ _3168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7944__A3 _3112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6948_ _1906_ _2071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5955__A2 _1119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6879_ _1973_ _2003_ _2004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_10_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8618_ _0063_ clknet_4_7_0_Clock B\[3\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6904__A1 _3510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8549_ _3737_ _3739_ _3740_ _0147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5891__A1 _3625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8582__CLK clknet_4_4_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6981__I _2102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8188__A3 _3002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7148__A1 _1530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7148__B2 _4069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7699__A2 _2851_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4676__I _3964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7623__A2 net34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7920_ _3031_ _3035_ _3086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6891__I _2014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7851_ _0479_ _0480_ _1732_ _1734_ _2867_ _3013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_64_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6802_ _1928_ _1929_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7782_ _0922_ _0923_ _1897_ _1898_ _3991_ _2940_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_4994_ _3979_ _0179_ _0180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6733_ _1863_ _1864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7139__A1 _4035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6664_ _1767_ _1798_ _1799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_109_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8403_ _3603_ _3605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5615_ _0759_ _0788_ _0789_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4360__B _3100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6595_ _3037_ _1731_ A\[0\]\[1\] _1732_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__4373__A1 _2745_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8334_ _3495_ _3508_ _3532_ _3533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5546_ _0663_ _0715_ _0722_ _0723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_121_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8265_ _3397_ _3404_ _3459_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5477_ _4071_ _0571_ _0654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7216_ _2268_ _2285_ _2345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4428_ _3718_ _3744_ _3745_ _3750_ _3751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_8196_ _3373_ _3383_ _3384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5873__A1 _4160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7147_ _2269_ _2270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4359_ _2856_ _3100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_101_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7078_ _2196_ _2197_ _2198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5625__A1 _4198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6029_ _1138_ _1191_ _1192_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_46_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5210__I _0390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4364__A1 _2971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5561__B1 _0539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5313__B1 _0036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7853__A2 _0388_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4667__A2 _3827_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5864__A1 _1028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4496__I _2982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5616__A1 _0773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7369__A1 _2440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6216__I _3972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8030__A2 _2350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5919__A2 _0723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6592__A2 _0000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4355__A1 _3037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5400_ _0576_ _0577_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6380_ _1372_ _1528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5698__A4 _0462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5331_ _0479_ _0480_ _3990_ _0508_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_55_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8097__A2 _3186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8050_ _0456_ C\[0\]\[8\] _3226_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5262_ _2695_ _0319_ _0440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7844__A2 _3005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6647__A3 _1723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4658__A2 _3780_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7001_ _2119_ _2121_ _2122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5855__A1 _4001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5193_ _2706_ _0374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5607__A1 _0309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7903_ _2981_ _3003_ _3068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4355__B A\[3\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7834_ _2942_ _2943_ _2995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8021__A2 _3179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5030__I _0025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7765_ _2861_ _2886_ _2922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4977_ _0149_ _0151_ _0163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7780__A1 _0391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6716_ _1706_ _1848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4594__B2 _3755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7696_ _0903_ _1811_ _2849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6647_ _0457_ C\[1\]\[2\] _1723_ _1781_ _1782_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__6335__A2 _0039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6578_ _0040_ _1716_ _1717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8317_ _3473_ _3476_ _3515_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5529_ _0703_ _0704_ _0705_ _0706_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_3_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6099__A1 _1245_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7835__A2 _2943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8248_ _3373_ _3383_ _3440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5846__A1 _4167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8179_ _3363_ _3292_ _3365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5205__I _3956_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8663__D _0118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7063__A3 _2050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6271__A1 _3883_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8620__CLK clknet_4_1_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7771__A1 _4158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4585__A1 _3902_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7523__A1 _2570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6877__A3 _2001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4888__A2 _4203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7826__A2 _2014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5301__A3 _0330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6655__B _3759_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7054__A3 _1807_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8251__A2 _1931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4900_ _4214_ _4215_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5880_ _0975_ _0977_ _1045_ _1046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_61_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6014__A1 _1029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4831_ _4065_ _4147_ _4148_ _4149_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_60_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6565__A2 _1704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7550_ _2661_ _2670_ _2703_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4762_ _4076_ _0020_ _4082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6501_ _1585_ _1588_ _1583_ _1645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7481_ _2627_ _2628_ _2629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_105_1144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4693_ _4013_ _3769_ _3967_ _3770_ _4014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4328__A1 _2745_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6432_ _1569_ _1577_ _1578_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_128_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6363_ _1418_ _1423_ _1512_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8102_ _3201_ _3279_ _3280_ _3281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5314_ _0489_ _4207_ _0378_ _0036_ _0491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6294_ _1429_ _1444_ _1445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_130_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5828__A1 _4139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8033_ _3201_ _3203_ _3206_ _3208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5245_ _0420_ _0421_ _0424_ _0425_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__8490__A2 _3669_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8643__CLK clknet_4_8_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5176_ _0342_ _0345_ _0355_ _0356_ _0357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4500__B2 _3788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6253__A1 _1400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4803__A2 _4100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6005__A1 _1028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7817_ _2924_ _2960_ _2976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7748_ _2848_ _2852_ _2903_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7679_ _2793_ _2832_ _2833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__4319__A1 _2545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6859__A3 _1980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8658__D _0127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8481__A2 _3666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7036__A3 _2156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7992__A1 _0050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_1_0_Clock_I clknet_3_0_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5819__B _0984_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7744__A1 _2846_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5770__A3 _0920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8568__D _0013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8666__CLK clknet_4_15_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5030_ _0025_ _0214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5038__A2 _0220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6981_ _2102_ _2103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4797__A1 _3846_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5932_ _1095_ _0713_ _0714_ _1097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_98_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8651_ _0093_ clknet_4_11_0_Clock C\[1\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5863_ _3777_ _3789_ _4182_ _1027_ _3926_ _1029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__6538__A2 _1679_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7735__A1 _2842_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7602_ _0223_ _0225_ _2754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_107_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4814_ _4128_ _4129_ _4131_ _4132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_37_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8582_ _0027_ clknet_4_4_0_Clock A\[3\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5794_ _0864_ _0865_ _0963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_72_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7533_ _2641_ _2643_ _2640_ _2686_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4745_ _3821_ _4066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7464_ _2561_ _2563_ _2612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4676_ _3964_ _3997_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8160__A1 _3261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6415_ _0327_ _1357_ _1358_ _1471_ _1351_ _1561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__4859__I _4092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7395_ _2476_ _2518_ _2537_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6710__A2 C\[1\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput18 net18 Result[11] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_116_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput29 net29 Result[6] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_6346_ _1493_ _1495_ _1496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_115_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6277_ _1426_ _1329_ _1427_ _1428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8463__A2 _3796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5277__A2 _0405_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8016_ _3947_ _0325_ _1755_ _3189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_131_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5228_ _0408_ _0409_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4808__B _4064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5159_ _0207_ _0324_ _0327_ _0329_ _0334_ _0339_ _0340_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai33_1
XFILLER_56_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8215__A2 _3404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6226__A1 _4173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4788__A1 _0056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5985__B1 _3625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7726__A1 _0775_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5201__A2 _0381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8689__CLK clknet_4_5_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4960__A1 _3809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4769__I _3542_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6701__A2 C\[1\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5268__A2 _0445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8206__A2 _1975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7965__A1 _3081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6768__A2 _1777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5440__A2 _0423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7717__A1 _2826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6940__A2 _1976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4530_ _2481_ _3853_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4951__A1 _4263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4461_ _3783_ _3784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6200_ _1242_ _1266_ _1355_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7180_ _2219_ _2288_ _2305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4392_ _2503_ _3456_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6131_ _1162_ _1189_ _1290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6456__A1 _1596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6062_ _1216_ _1223_ _1224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_113_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5013_ _3133_ _0199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6759__A2 _1853_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6964_ _2086_ _2087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5431__A2 _0607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5915_ _1056_ _1078_ _1079_ _1080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_34_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6895_ _1942_ _2006_ _2018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7708__A1 _0751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5846_ _4167_ _4187_ _1012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8634_ _0108_ clknet_4_11_0_Clock C\[0\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7184__A2 _2242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5777_ _0024_ _0048_ _0946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8565_ _0010_ clknet_4_0_0_Clock A\[1\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7516_ C\[1\]\[14\] _0186_ _2667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4728_ _3959_ _3963_ _4049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8496_ _3694_ _3695_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7447_ _2535_ _2593_ _2594_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_68_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4659_ _3980_ _3981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6695__A1 _4215_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7378_ _2476_ _2518_ _2519_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_66_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6329_ _1374_ _1479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5670__A2 _0498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7947__A1 _3019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8524__I _3683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8671__D _0065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7411__A3 _2552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8372__A1 _3446_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8372__B2 _3498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7714__A4 _0002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6979__I _2100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5186__A1 _3845_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8124__A1 _0487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4499__I _3821_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6219__I _1247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4464__A3 _3748_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7938__A1 _0481_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7938__B2 _0382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8581__D _0026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5700_ _3876_ _0462_ _0842_ _0795_ _0873_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_108_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6680_ _0202_ _0010_ _1812_ _3510_ _1813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_52_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8363__A1 _3555_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5631_ _0471_ _0483_ _0455_ _0805_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_73_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6913__A2 _2014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8350_ _3547_ _3548_ _3549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5562_ _0512_ _4015_ _0537_ _0533_ _0739_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__8115__A1 _3278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7301_ _3971_ C\[1\]\[10\] _2155_ _2185_ _2436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4513_ _3826_ _3834_ _3836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8281_ _3474_ _3475_ _3476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5493_ _0622_ _0669_ _0670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_89_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7232_ _2359_ _2360_ _2361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4444_ _3766_ _3767_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_144_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7163_ _2245_ _2248_ _2286_ _2288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_63_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4375_ _3260_ _3271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_63_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6114_ _1272_ _1273_ _1274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7094_ _2207_ _2213_ _2214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_100_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6045_ _1055_ _1063_ _1207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5652__A2 _0033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7929__A1 _0577_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7996_ _3158_ _3160_ _3166_ _3167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_1607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5404__A2 _0573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6947_ _1991_ _1993_ _2000_ _2070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4612__B1 _3829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6878_ _1974_ _1976_ _2002_ _2003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__7157__A2 _2151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8617_ _0062_ clknet_4_9_0_Clock B\[3\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5829_ _4132_ _4143_ _0995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6904__A2 _0013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8548_ _0107_ _3714_ _3740_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8106__A1 _3283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8479_ _3673_ _3679_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7865__B1 _1781_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7851__C _2867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8666__D _0121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5340__A1 _0512_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8409__A2 _3566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5340__B2 _3976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5891__A2 _0750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7093__A1 _2211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6840__A1 _2460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_78 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8345__A1 _3492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7148__A2 _1826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5159__A1 _0207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5159__B2 _0334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6659__A1 _1727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8576__D _0021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5331__A1 _0479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5882__A2 _4260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7084__A1 _3889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4692__I A\[2\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7850_ _2949_ _3010_ _3011_ _2957_ _2945_ _3012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_63_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7387__A2 _2455_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6801_ _1927_ _1928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5398__A1 _0574_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7781_ _0348_ _0352_ _1847_ _1850_ _3593_ _2939_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_17_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4993_ B\[1\]\[0\] _3764_ _3391_ _3765_ _0179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_90_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6732_ _1862_ _1863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__8336__A1 _3492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7139__A2 _1746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6663_ _1774_ _1797_ _1798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5614_ _0785_ _0787_ _0788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6898__A1 _1944_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8402_ _3598_ _3602_ _3603_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6594_ _1709_ _1731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_34_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8333_ _3512_ _3530_ _3532_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4373__A2 _3048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5545_ _0717_ _0719_ _0721_ _0722_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_117_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8264_ _3407_ _3408_ _3457_ _3458_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5476_ _0650_ _0652_ _0653_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5322__A1 _0419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7215_ _2268_ _2285_ _2344_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4427_ _3749_ _3750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8195_ _3377_ _3382_ _3383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_87_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7146_ _4001_ _1319_ _1980_ _1999_ _2269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_101_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4358_ _3067_ _3078_ _2631_ _3089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_99_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7077_ _2116_ _2129_ _2197_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8275__S _3469_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4289_ net2 _2362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_58_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5625__A2 _0462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6028_ _1140_ _1190_ _1191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_58_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5389__A1 _0564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7979_ _3148_ _0963_ _3149_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8327__A1 _0038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7418__I _2163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4364__A2 _3144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5561__A1 _0512_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5561__B2 _4015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5313__A1 _4207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5313__B2 _0489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5864__A2 _1029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7369__A2 _2441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4355__A2 _3048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5552__A1 _0636_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5330_ _3813_ _0506_ _0507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5261_ _0407_ _0438_ _0439_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5304__A1 _3997_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6647__A4 _1781_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7000_ _4113_ _2120_ _2048_ _2121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5855__A2 _3948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5192_ _0341_ _0371_ _0372_ _0373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7902_ _2994_ _3007_ _3065_ _3066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5311__I _0488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7833_ _2926_ _2931_ _2994_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7764_ _2909_ _2920_ _2921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4976_ _0152_ _0153_ _0162_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_11_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7780__A2 _0400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6715_ _1846_ _1847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4594__A2 _3753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8572__CLK clknet_4_3_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7695_ _2770_ _2777_ _2813_ _2848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_109_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6646_ _1780_ _1781_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__7532__A2 _2592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6577_ _1715_ _1716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8316_ _3465_ _3472_ _3514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5528_ _4015_ _0393_ _0705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7296__A1 _2364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8247_ _3377_ _3382_ _3439_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5459_ _0634_ _0572_ _0635_ _0636_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5846__A2 _4187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8178_ _3363_ _3292_ _3364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7129_ _1899_ _2250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6271__A2 _3899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8548__A1 _0107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_3_1_0_Clock_I clknet_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7220__A1 _4035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7771__A2 _0751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5782__A1 _0016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7523__A2 _2604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6731__B1 _1698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7039__A1 _4003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6227__I _0718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8595__CLK clknet_4_0_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7211__A1 _2334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8442__I _3645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4830_ _4050_ _4099_ _4148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5773__A1 _0937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4761_ _4081_ _0020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6500_ _1642_ _1643_ _1644_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7480_ _1530_ _0006_ _2628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_14_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4692_ A\[2\]\[6\] _4013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4328__A2 _2755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5525__A1 _3922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6431_ _1575_ _1576_ _1577_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_105_1178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6362_ _1425_ _1446_ _1510_ _1511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5313_ _4207_ _0378_ _0036_ _0489_ _0490_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8101_ _3203_ _3206_ _3280_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6293_ _1433_ _1443_ _1444_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_143_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5828__A2 _4142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8032_ _3204_ _3205_ _3206_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5244_ _0422_ _0423_ _0424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4500__A2 _3787_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5175_ _3773_ _0356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6253__A2 _1404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7450__A1 _2573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7202__A1 _4195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6005__A2 _1029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8352__I _2665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7816_ _2924_ _2960_ _2975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7753__A2 _2811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7747_ _2848_ _2852_ _2902_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4959_ _3953_ _4273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7678_ _2762_ _2796_ _2831_ _2832_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_138_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6629_ _0211_ _0009_ _1763_ _1764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6859__A4 _1983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7269__A1 _4133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5216__I _3840_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8674__D _0081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7036__A4 _1826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6795__A3 _1922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7992__A2 _0013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5204__B1 _0384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4558__A2 _3879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_5_0_Clock_I clknet_3_2_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5126__I _0307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8584__D _0029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7432__A1 _3883_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6980_ _2101_ _2102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6786__A3 _0011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5931_ _0713_ _0714_ _1095_ _1096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4797__A2 _4028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8650_ _0092_ clknet_4_11_0_Clock C\[1\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5862_ _3777_ _3789_ _4182_ _1027_ _1028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_90_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7601_ _2753_ _0069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4813_ _3849_ _4130_ _4131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8581_ _0026_ clknet_4_4_0_Clock A\[3\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5793_ _0918_ _0960_ _0961_ _0962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7532_ _2588_ _2592_ _2683_ _2684_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4744_ _4053_ _4055_ _4064_ _4065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_124_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7463_ _2550_ _2608_ _2609_ _2558_ _2566_ _2611_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_4675_ _3989_ _3833_ _3995_ _3996_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6414_ _1559_ _1498_ _1560_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8610__CLK clknet_4_11_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7394_ _2411_ _2473_ _2536_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_66_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput19 net19 Result[12] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_6345_ _1360_ _1385_ _1494_ _1495_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4721__A2 _3987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5036__I _3882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6276_ _1315_ _1328_ _1427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_131_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8015_ _2998_ _3186_ _3187_ _3095_ _3188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5227_ _0307_ _0408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7671__A1 _1479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7251__I _2381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5158_ _0022_ _0339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6226__A2 _0039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5089_ _0270_ _0271_ _0272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_16_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4788__A2 _4107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5985__A1 _4195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5985__B2 _4202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7726__A2 _1783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8669__D _0124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4960__A2 _4273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6701__A3 _1723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7662__A1 _0348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7414__A1 _2550_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7965__A2 _3135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7717__A2 _1848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5728__A1 _0774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8633__CLK clknet_4_11_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8579__D _0024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4951__A2 _4264_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4460_ _2352_ _3748_ _3782_ _3783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_116_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5900__A1 _0689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4391_ _2276_ _3445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_125_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6130_ _1162_ _1189_ _1289_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6061_ _1221_ _1222_ _1223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7653__A1 _0897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5012_ _0192_ _0196_ _0197_ _0198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6963_ _1981_ _1982_ _3990_ _2086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8702_ _0148_ clknet_4_13_0_Clock net22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5914_ _3897_ _0051_ _1079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6894_ _1942_ _2006_ _2017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7708__A2 _1746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8633_ _0107_ clknet_4_11_0_Clock C\[0\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5845_ _0996_ _1010_ _1011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8564_ _0009_ clknet_4_1_0_Clock A\[1\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6392__A1 _1538_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5776_ _0945_ _0048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7515_ _1597_ C\[1\]\[14\] B\[1\]\[7\] _2665_ _2666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4727_ _3932_ _4044_ _4046_ _4047_ _3963_ _4048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_8495_ _3673_ _3674_ _3694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7446_ _2588_ _2592_ _2593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4658_ B\[1\]\[6\] _3780_ _3572_ _3783_ _3980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__6695__A2 _0001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7377_ _2490_ _2517_ _2518_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4589_ _3682_ _3909_ _3910_ _3911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6328_ _3636_ _0711_ _1478_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6259_ _1167_ _1188_ _1411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_88_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7947__A2 _1980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8656__CLK clknet_4_6_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6383__A1 _4070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5186__A2 _0362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8124__A2 _1986_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8507__S0 _3704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4464__A4 _3782_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7938__A2 _1841_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5630_ _0791_ _0798_ _0803_ _0804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5177__A2 _2578_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5561_ _0512_ _0537_ _0539_ _4015_ _0738_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7300_ _0473_ C\[1\]\[10\] _3974_ _2435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6126__A1 _1145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4512_ _3826_ _3834_ _3835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5492_ _0625_ _0668_ _0669_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8280_ _0384_ _2501_ _3475_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7231_ _1319_ _1791_ _1983_ _1163_ _2360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_89_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4443_ _3763_ _3764_ _3196_ _3765_ _3766_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_4374_ _2805_ net10 _3260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7162_ _2264_ _2268_ _2285_ _2286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_98_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6113_ _1205_ _1206_ _1271_ _1273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_112_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7093_ _2211_ _2212_ _2213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6044_ _1051_ _1115_ _1206_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8679__CLK clknet_4_7_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7929__A2 _1823_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4860__A1 _3978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8051__A1 _3926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7995_ _3164_ _3165_ _3166_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_93_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6946_ _1991_ _1993_ _2000_ _2069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_82_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4612__B2 _3756_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6877_ _1979_ _1989_ _2001_ _2002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_126_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8616_ _0061_ clknet_4_1_0_Clock B\[3\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5828_ _4139_ _4142_ _0994_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6365__A1 _3900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8547_ _3693_ _3738_ _3708_ _3739_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5759_ _0906_ _0907_ _0902_ _0929_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_124_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8478_ _3667_ _3678_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_11_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7865__A1 _0720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7429_ _2559_ _2574_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7865__B2 _0383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4679__A1 _3997_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5340__A2 _0466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7617__A1 _0897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8290__A1 _3424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8682__D _0075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6840__A2 _1811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5159__A2 _0324_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5159__B3 _0339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4906__A2 _4220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6659__A2 _1729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5331__A2 _0480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7084__A2 _2203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8592__D _0037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6831__A2 _1912_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4842__A1 _4157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8033__A1 _3201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6800_ _1926_ _3775_ _1861_ _1698_ _3829_ _1927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_91_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6595__A1 _3037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7780_ _0391_ _0400_ _1713_ _1735_ _2938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_91_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4992_ _0176_ _0177_ _0178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6731_ _1860_ _2674_ _1861_ _1698_ _3802_ _1862_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_90_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6662_ _1793_ _1796_ _1797_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_108_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8401_ _3599_ _3600_ _3601_ _3602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5613_ _0329_ _0786_ _0787_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_20_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6593_ _1727_ _1729_ _1730_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5309__I _0400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8332_ _3513_ _3529_ _3530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_30_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5544_ _4169_ _0720_ _0721_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8263_ _3406_ _3409_ _3457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5475_ _3772_ _0569_ _0651_ _3956_ _0652_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_144_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7214_ _2325_ _2342_ _2343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4426_ _3746_ _3748_ _2567_ _3749_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5322__A2 _0498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8194_ _3379_ _3381_ _3382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_63_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7145_ _2154_ _2266_ _2267_ _2268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4357_ _2805_ net6 _3078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_86_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8272__A1 _0457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7076_ _2118_ _2128_ _2196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4288_ _2254_ _2352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_115_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6027_ _1160_ _1162_ _1189_ _1190_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_39_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5389__A2 _0565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7978_ _0893_ _0962_ _3148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6586__A1 _3759_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6929_ _4133_ _1882_ _2052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8327__A2 _3302_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5010__A1 _0193_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5561__A2 _0537_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8677__D _0084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7838__A1 _2236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5313__A2 _0378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7066__A2 _2184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4793__I _4112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5129__I _0303_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7829__A1 _2979_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8587__D _0032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5260_ _4262_ _0051_ _0438_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5304__A2 _0481_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5191_ _0366_ _0370_ _0372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8006__A1 _3126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7901_ _2997_ _3006_ _3065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7832_ _2933_ _2959_ _2991_ _2992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7763_ _2910_ _2918_ _2920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4975_ _4269_ _0160_ _0161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8309__A2 _3505_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5240__A1 _0419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6714_ _2492_ _1731_ A\[0\]\[3\] _1846_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7780__A3 _1713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7694_ _0945_ _0011_ _2797_ _2847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_123_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6645_ _1779_ _1780_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6576_ _1714_ _1715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6740__A1 _1760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4878__I _2963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8315_ _3474_ _3475_ _3513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_117_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5527_ _4010_ _0401_ _0704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8493__A1 _3683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8246_ _3436_ _3437_ _3438_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7296__A2 _2368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5458_ _3965_ _4213_ _0632_ _0633_ _0635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_133_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4409_ _3625_ _3636_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8177_ _3289_ _3363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5389_ _0564_ _0565_ _0566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_8_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7128_ _4076_ _0004_ _2141_ _2249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7048__A2 _2158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5059__A1 _4113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7059_ _2179_ _1823_ _1998_ _3785_ _2180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_101_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8548__A2 _3714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6559__A1 _2481_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7220__A2 _1757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7771__A3 _2237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_5_0_Clock_I clknet_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5782__A2 _0757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6731__A1 _1860_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6731__B2 _3802_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8484__A1 _3683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7039__A2 _1791_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6952__B A\[0\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4760_ _3778_ _4080_ _4081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5773__A2 _0181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4691_ _3832_ _4012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8172__B1 _3284_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6430_ _1375_ _1482_ _1484_ _1487_ _1576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6722__A1 _1836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4328__A3 _2764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5525__A2 _3772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6361_ _1428_ _1445_ _1510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_127_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8100_ _3203_ _3206_ _3279_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5312_ _3922_ _0489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6292_ _1434_ _1442_ _1443_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_115_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8031_ _0924_ _2404_ _3205_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5243_ _0360_ _0423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8227__A1 _3354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5174_ _0354_ _0355_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6789__A1 _4113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5461__A1 _3805_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7815_ _2972_ _2973_ _2974_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5213__A1 _0386_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7746_ _2799_ _2899_ _2900_ _2901_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5764__A2 _0919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6961__A1 _3998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4958_ _4270_ _4271_ _4272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_123_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7677_ _2802_ _2806_ _2830_ _2831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_4889_ _4199_ _4204_ _4205_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6628_ _0208_ _1759_ _1763_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_140_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6559_ _2481_ _3746_ _3747_ _2287_ _1699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_134_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7269__A2 _1864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8229_ _3348_ _3419_ _3420_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_12_0_Clock_I clknet_3_6_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8218__A1 _0488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5232__I _0362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7992__A3 _3093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5204__A1 _0374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5204__B2 _3997_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6952__A1 _2745_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_9_0_Clock_I clknet_3_4_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6180__A2 _1197_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4311__I _2589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8209__A1 _1178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5691__A1 _0835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8562__CLK clknet_4_10_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7432__A2 _2126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5930_ _3876_ _1094_ _0662_ _1095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_18_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5861_ _0513_ C\[3\]\[9\] _1027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7196__A1 _2234_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7600_ _2741_ _2752_ _2753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4812_ _3293_ _4130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8580_ _0025_ clknet_4_1_0_Clock A\[3\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5792_ _0888_ _0891_ _0961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6943__A1 _3818_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7531_ _2641_ _2643_ _2640_ _2683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4743_ _4057_ _4058_ _4063_ _4064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_30_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7462_ _2551_ _2557_ _2609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4674_ _3800_ _0042_ _3806_ _3995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_135_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6413_ _1464_ _1559_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7393_ _2529_ _2533_ _2535_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6344_ _1361_ _1362_ _1384_ _1494_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8448__A1 _1688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6275_ _1311_ _1426_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8014_ _1184_ _0326_ _2911_ _1701_ _0577_ _3187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_5226_ _3848_ _0320_ _0407_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4377__B _3100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5157_ _0338_ _0022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5088_ _4266_ _4267_ _0271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4891__I _3840_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5985__A2 _3897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7187__A1 _3026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6934__A1 _2051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7729_ _2880_ _2884_ _2885_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_90_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6611__I _1747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5227__I _0307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6701__A4 _0000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8439__A1 _3627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8585__CLK clknet_4_6_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7111__A1 _2184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7662__A2 _0352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5425__A1 _0536_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5976__A2 _0989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7178__A1 _2205_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6925__A1 _2031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5728__A2 _0899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4390_ _3423_ _3434_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8595__D _0040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7102__A1 _2178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6060_ _1219_ _1220_ _1222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7653__A2 _1704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5664__A1 _0833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input8_I X[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5011_ _0183_ _0187_ _0197_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6962_ _2082_ _2084_ _2085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5600__I _3964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8701_ _0147_ clknet_4_13_0_Clock net21 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5913_ _4026_ _0409_ _1078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6893_ _1934_ _2008_ _2015_ _2016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_22_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8632_ _0106_ clknet_4_11_0_Clock C\[0\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5844_ _0998_ _1009_ _1010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5719__A2 _0891_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6916__A1 _2028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8563_ _0008_ clknet_4_0_0_Clock A\[1\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5775_ _0467_ _0945_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6392__A2 _0023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7514_ _2501_ _2665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4726_ _3993_ _4002_ _3950_ _4047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_8494_ _3692_ _3693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7445_ _2467_ _2590_ _2591_ _2592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_68_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4657_ _3978_ _3979_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7376_ _2493_ _2516_ _2517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4588_ _3887_ _3908_ _3910_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4886__I _3844_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6327_ _1366_ _1376_ _1476_ _1477_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6258_ _1294_ _1304_ _1410_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5655__A1 _3875_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5209_ _3701_ _0389_ _0390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6189_ _1225_ _1344_ _1345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5510__I _0444_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6383__A2 _1530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7580__A1 _1598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4394__A1 _3434_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8507__S1 _3679_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8268__I _0632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5646__A1 _0587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6071__A1 _3898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8600__CLK clknet_4_9_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5177__A3 _0346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4385__A1 _3358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5560_ _4061_ _0539_ _0737_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4511_ _3758_ _3827_ _3833_ _3834_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5491_ _0641_ _0645_ _0667_ _0668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_129_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7230_ _1985_ _1529_ _1975_ _2087_ _2359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4442_ _3755_ _3765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__7874__A2 _3012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7161_ _2272_ _2284_ _2285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_113_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4373_ _2745_ _3048_ _2534_ A\[3\]\[5\] _3249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_98_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6112_ _1205_ _1206_ _1271_ _1272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7626__A2 _2777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7092_ _3240_ _2126_ _2212_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6043_ _1053_ _1114_ _1205_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4860__A2 _4091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7994_ _0049_ _2203_ _3165_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6945_ _1984_ _2067_ _2068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_81_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4612__A2 _3754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6876_ _1905_ _1994_ _2000_ _2001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5827_ _4149_ _0989_ _0990_ _0991_ _0992_ _0993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_50_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8615_ _0060_ clknet_4_1_0_Clock B\[3\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6365__A2 _1419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8546_ _0122_ _0077_ _3695_ _3738_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5758_ _0016_ _0925_ _0927_ _0928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_72_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4709_ _4027_ _4029_ _4030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8477_ _0124_ _3669_ _3671_ _3676_ _3677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7314__A1 _2387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5689_ _0856_ _0860_ _0861_ _0862_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_68_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7428_ _2571_ _2572_ _2573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7865__A2 _2771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4679__A2 _3825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7359_ _2496_ _2497_ _2498_ _2499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7617__A2 _1703_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8623__CLK clknet_4_0_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8042__A2 _3210_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5800__A1 _0821_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5159__A3 _0327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7305__A1 _4085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7856__A2 _0505_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5867__A1 _1024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5619__A1 _3973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8281__A2 _3475_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4842__A2 _4159_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6044__A1 _1051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4991_ _4232_ _4258_ _0177_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6595__A2 _1731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7792__A1 _0383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6730_ _1699_ _1861_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_90_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6661_ _1719_ _1794_ _1795_ _1796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5612_ _0022_ _0436_ _0786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8400_ _3462_ _2665_ _3601_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6592_ _4157_ _0000_ _1728_ _1729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_121_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8331_ _3516_ _3528_ _3529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5543_ _0571_ _0720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8262_ _3390_ _3453_ _3454_ _3455_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5474_ _0648_ _0651_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7213_ _2327_ _2340_ _2342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4425_ _3747_ _3748_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
X_8193_ _0408_ _1929_ _3381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5322__A3 _0464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7144_ _2158_ _2166_ _2167_ _2267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8646__CLK clknet_4_8_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4356_ _2786_ _3067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7075_ _2195_ _0099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4287_ _2330_ net7 _2341_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_140_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6283__A1 _0045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6026_ _1167_ _1188_ _1189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7977_ _3147_ _0084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6928_ _3793_ _3861_ _2050_ _2051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_126_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6859_ _4001_ _4150_ _1980_ _1983_ _1984_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__7535__A1 _2646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4349__A1 _2982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4349__B2 B\[3\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8529_ _0116_ _3723_ _3714_ _3724_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7838__A2 _0307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5235__I _0415_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8693__D _0139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8015__A2 _3186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6026__A1 _1167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7774__A1 _2926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4314__I _2621_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5001__A2 _0186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8669__CLK clknet_4_15_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4760__A1 _3778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5145__I _0326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4512__A1 _3826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5190_ _0366_ _0370_ _0371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8254__A2 _3446_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6265__A1 _0061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5068__A2 _0249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7900_ _2985_ _2986_ _3063_ _3064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6017__A1 _4045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7831_ _2934_ _2990_ _2958_ _2991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7765__A1 _2861_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4579__A1 _3889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4974_ _0154_ _0156_ _0160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7762_ _2916_ _2917_ _2918_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_51_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5240__A2 _0414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6713_ _1843_ _1844_ _1845_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7693_ _2798_ _2801_ _2843_ _2844_ _2846_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__7517__A1 _1533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6644_ _1776_ _1778_ _3760_ _1779_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6575_ _1713_ _1714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8314_ _3458_ _3509_ _3511_ _3512_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5526_ _0652_ _0654_ _0702_ _0703_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8245_ _3386_ _3414_ _3437_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5457_ _3965_ _0632_ _0633_ _4213_ _0634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_133_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4408_ _3615_ _3625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4503__A1 _3814_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8176_ _3296_ _3360_ _3361_ _3362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5388_ _2755_ _3893_ _0380_ _0565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_120_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7127_ _2055_ _0004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4339_ _2878_ _2889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5059__A2 _0200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7058_ _3866_ _2179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4806__A2 _4037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6009_ _4172_ _4062_ _1172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6008__A1 _1024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6559__A2 _3746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7756__A1 _4158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8181__A1 _0899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8688__D _0134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6731__A2 _2674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4742__A1 _4012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8484__A2 _3674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7039__A3 _2159_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5773__A3 _0920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4690_ _3952_ _4009_ _4010_ _4011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8172__A1 _0897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8598__D _0043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6722__A2 _1853_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6360_ _1416_ _1424_ _1509_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4733__A1 _3825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5311_ _0488_ _0036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8475__A2 _3674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6291_ _1436_ _1440_ _1441_ _1442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_143_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8030_ _0822_ _2350_ _3204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5242_ _3831_ _0422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4497__B1 _3819_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5173_ _0353_ _0354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6789__A2 _1762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7986__A1 _0049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput1 Enable net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_84_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5461__A2 _0487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7814_ _2909_ _2920_ _2973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5213__A2 _0393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7745_ _2846_ _2890_ _2900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4957_ _3814_ _4007_ _4271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8538__I0 _0120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5764__A3 _0932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6961__A2 _1781_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7676_ _2808_ _2814_ _2829_ _2830_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_4888_ _4201_ _4203_ _4204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_137_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6627_ _1762_ _0009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6558_ _3779_ _3445_ _3782_ _1698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_106_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5509_ _0608_ _0610_ _0685_ _0686_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6489_ _1573_ _1574_ _1633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6477__A1 _1619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8228_ _3351_ _3418_ _3419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_133_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8218__A2 _3302_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8159_ _3339_ _3332_ _3342_ _3343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_86_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5204__A2 _0378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8529__I0 _0116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6952__A2 _1777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4799__I _4116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7901__A1 _2997_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4715__A1 _4033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6963__B _3990_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5860_ _4183_ _4185_ _1025_ _1026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4811_ _4112_ _3604_ _4129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5791_ _0934_ _0958_ _0959_ _0960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6943__A2 _1907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7530_ _2650_ _2681_ _2682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4742_ _4012_ _4062_ _4063_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8145__A1 _3274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7461_ _2551_ _2557_ _2608_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4673_ _3994_ _0042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6412_ _1468_ _1497_ _1558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4706__A1 _2449_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7392_ _2523_ _2531_ _2532_ _2533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6343_ _1490_ _1492_ _1493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_66_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6274_ _1416_ _1424_ _1425_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_131_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5225_ _0396_ _0405_ _0406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8013_ _3947_ _0576_ _2050_ _3186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__5131__A1 _2599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5156_ _0336_ _0337_ _0338_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7959__A1 _0434_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5087_ _0239_ _0243_ _0270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6631__A1 _4116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_13_0_Clock clknet_3_6_0_Clock clknet_4_13_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_53_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7187__A2 _1929_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5989_ _4141_ _1150_ _1151_ _1005_ _1152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XPHY_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7728_ _2881_ _2882_ _2883_ _2884_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_7659_ _0752_ _1703_ _1747_ _0896_ _2812_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_14_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5370__A1 _0492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5243__I _0360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5425__A2 _0543_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8503__B _3700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6802__I _1928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8127__A1 _3228_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5361__A1 _4130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5153__I _3778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ _0193_ _0194_ _0195_ _0196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__5664__A2 _0834_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8464__I net14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6961_ _3998_ _1781_ _2083_ _2084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8700_ _0146_ clknet_4_13_0_Clock net20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5912_ _0701_ _0706_ _1076_ _1077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6892_ _1937_ _2007_ _2015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8631_ _0105_ clknet_4_10_0_Clock C\[0\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5843_ _1001_ _1008_ _1009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_50_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8562_ _0007_ clknet_4_10_0_Clock A\[0\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5774_ _0939_ _0943_ _0944_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7029__B A\[0\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7513_ _2626_ _2662_ _2664_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4725_ _3820_ _4045_ _3937_ _4046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_8493_ _3683_ _3667_ _3692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7444_ _2469_ _2520_ _2591_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4656_ _3812_ _3978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4587_ _3887_ _3908_ _3909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_66_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7375_ _2507_ _2515_ _2516_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_131_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6326_ _1378_ _1382_ _1476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_115_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6159__I _1164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6257_ _1288_ _1407_ _1408_ _1409_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5655__A2 _0364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5208_ _0387_ _0388_ _0389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_88_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6188_ _1269_ _1344_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5139_ _3875_ _0320_ _0321_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6604__A1 _0211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4407__I _3604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8357__A1 _1528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6622__I _1757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8109__A1 _3088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7580__A2 C\[0\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4394__A2 _2352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5591__A1 _0356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5894__A2 _0734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4697__A3 _4017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7096__A1 _2135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6071__A2 _0607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8348__A1 _3512_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7020__A1 _3980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4909__A1 _4222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4385__A2 _3369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4510_ _3831_ _3832_ _3833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5490_ _0655_ _0666_ _0667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_89_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8520__A1 _0114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4441_ _3753_ _3764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_89_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7874__A3 _3038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7160_ _2274_ _2280_ _2283_ _2284_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_4372_ _3229_ _3240_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6111_ _1210_ _1213_ _1270_ _1271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_113_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7087__A1 _2174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7091_ _3004_ _1814_ _2208_ _2210_ _2211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7626__A3 _2778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6042_ _1204_ _0073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4860__A3 _4176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7993_ _3161_ _3162_ _3164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6944_ _2065_ _2066_ _2067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_82_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6875_ _3798_ _1999_ _2000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__8575__CLK clknet_4_1_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8614_ _0059_ clknet_4_3_0_Clock B\[3\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5826_ _4146_ _0992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8545_ _3719_ _0092_ _3737_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4376__A2 _3271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5757_ _0872_ _0874_ _0926_ _0927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_72_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4708_ _3846_ _4028_ _4029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8476_ _3675_ _3676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5688_ _0789_ _0810_ _0861_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8511__A1 _0098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7427_ _2410_ _2487_ _2572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8369__I _1094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4639_ _3960_ _3961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_135_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5876__A2 _1041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4679__A3 _3999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7358_ _4090_ C\[1\]\[11\] _2156_ _2164_ _2498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6309_ _1346_ _1387_ _1459_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_103_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7289_ _4034_ _1808_ _2423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6825__A1 _1948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6617__I _2867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8042__A3 _3214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8502__A1 _0095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7305__A2 _1962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4600__I _3921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8598__CLK clknet_4_9_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7241__A1 _2358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4990_ _0159_ _0174_ _0175_ _0176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_63_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6660_ _1727_ _1729_ _1737_ _1795_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_5611_ _0773_ _0783_ _0784_ _0785_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5555__A1 _3304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4358__A2 _3078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6591_ _1371_ C\[1\]\[1\] _0468_ _1728_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
X_8330_ _3517_ _3527_ _3528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_34_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5542_ _4218_ _0718_ _0719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8261_ _3394_ _3411_ _3454_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5473_ _0386_ _4273_ _0647_ _0649_ _0650_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_117_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4424_ _2265_ _3747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_8
X_7212_ _2332_ _2339_ _2340_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5858__A2 _1023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8192_ _3375_ _3378_ _3379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_99_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7143_ _2166_ _2167_ _2158_ _2266_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4355_ _3037_ _3048_ _2534_ A\[3\]\[1\] _3056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_119_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7074_ _2106_ _2110_ _2194_ _2195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_119_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4286_ _2319_ _2330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_115_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7042__B _3100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7480__A1 _1530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6283__A2 _1037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6025_ _1171_ _1187_ _1188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_45_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4294__A1 _2341_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6035__A2 _1197_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7232__A1 _2359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7976_ _0176_ _0177_ _3146_ _3147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_1407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5794__A1 _0864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6927_ _1744_ _2050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_70_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6858_ _1981_ _1982_ _1983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_50_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5809_ _4111_ _0973_ _0974_ _4119_ _4109_ _0975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__4349__A2 _2908_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6789_ _4113_ _1762_ _1824_ _1917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_13_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8528_ _3720_ _3722_ _3723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7299__A1 _1018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8459_ _3661_ _3799_ _0041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7838__A3 _2911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5849__A2 _4183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5482__B1 _0658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7774__A2 _2931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5537__A1 _4198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5537__B2 _0469_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4760__A2 _4080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4330__I _2786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5161__I _0310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7214__A1 _2325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6017__A2 _4067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7830_ _2879_ _2885_ _2990_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_97_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4579__A2 _3900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7761_ _2759_ _1931_ _2917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4973_ _4269_ _0157_ _0158_ _0159_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6712_ _4009_ _1841_ _1842_ _3975_ _1844_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4505__I A\[2\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7692_ _2806_ _2830_ _2844_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7517__A2 _2152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6643_ _3196_ _1777_ _1778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5528__A1 _4015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6574_ _1708_ _1712_ _1713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__8613__CLK clknet_4_1_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8313_ _3461_ _3477_ _3511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5525_ _3922_ _3772_ _0646_ _0651_ _0702_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_117_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5336__I _3854_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8244_ _3388_ _3412_ _3436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5456_ _0568_ _0633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4407_ _3604_ _3615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4503__A2 _3818_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5700__A1 _3876_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8175_ _3299_ _3327_ _3361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5387_ _3853_ _2578_ _0346_ B\[0\]\[7\] _0564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_87_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7126_ _2144_ _2246_ _2247_ _2248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4338_ _2775_ _2845_ _2867_ _2878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7057_ _2175_ _2176_ _2177_ _2178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_46_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6008_ _1024_ _1032_ _1170_ _1171_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7205__A1 _2179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6559__A3 _3747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7756__A2 _0761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7959_ _0434_ _2281_ _3129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_91_38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5519__A1 _0645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8181__A2 _2614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4742__A2 _4062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5690__B _0861_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6247__A2 _1197_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6805__I _1931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5758__A1 _0016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4325__I _2737_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4430__A1 _2737_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8636__CLK clknet_4_1_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8172__A2 _2390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5525__A4 _0651_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5930__A1 _3876_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5310_ _0487_ _0488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6290_ _0335_ _3981_ _0337_ _1441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_46_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5241_ _3806_ _0415_ _0421_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7371__I _2087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4497__A1 B\[1\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4497__B2 _3784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5172_ _0348_ _0352_ _3593_ _0353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_116_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6789__A3 _1824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7986__A2 _0014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput2 K[0] net2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_68_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7813_ _2910_ _2918_ _2972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5749__A1 _0336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7744_ _2846_ _2890_ _2899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_1272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4956_ _3762_ _3922_ _3767_ _4270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_127_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8538__I1 _0075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7675_ _2819_ _2823_ _2828_ _2829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_20_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4887_ _4070_ _4202_ _3856_ _3857_ _4203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_123_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6626_ _1761_ _1762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_119_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6557_ _1696_ _1697_ _0079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5508_ _0590_ _0609_ _0685_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_1519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6488_ _1570_ _1629_ _1631_ _1632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6477__A2 _1621_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8227_ _3354_ _3417_ _3418_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_79_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5439_ _4056_ _0354_ _0616_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4488__A1 _3758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8158_ _3334_ _3340_ _3341_ _3342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7109_ _2227_ _2228_ _2229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_75_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8089_ _0318_ _1928_ _3267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5988__A1 _2695_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5988__B2 _4031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8659__CLK clknet_4_7_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7729__A2 _2884_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output22_I net22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8699__D _0145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4963__A2 _4274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6165__A1 _0473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7901__A2 _3006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4715__A2 _4035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4479__A1 _2233_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7417__A1 _1295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8090__A1 _3092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8393__A2 _0015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4810_ _3841_ _3844_ _4128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5790_ _0867_ _0887_ _0916_ _0959_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_1590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4741_ _4061_ _4062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7460_ _2602_ _2606_ _2607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4672_ _3993_ _3786_ _3994_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6411_ _1557_ _0076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4706__A2 _4026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7391_ _2465_ _2530_ _2521_ _2532_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6342_ _1369_ _1476_ _1491_ _1383_ _1365_ _1492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__6459__A2 _1540_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6273_ _1418_ _1423_ _1424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_115_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8012_ _3180_ _3183_ _3184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_102_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5224_ _0399_ _0402_ _0404_ _0405_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_29_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7408__A1 _1530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5155_ A\[2\]\[6\] _4078_ net44 _4077_ _0337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_99_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7959__A2 _2281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5086_ _0268_ _0165_ _0162_ _0269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__6631__A2 _1703_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8384__A2 _3538_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5198__A2 _2578_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5988_ _2695_ _3872_ _4137_ _4031_ _1151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6934__A3 _2056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7727_ C\[0\]\[4\] _4239_ _2883_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4939_ _4252_ _4253_ _4254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8136__A2 _3311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7658_ _0050_ _1762_ _2810_ _2811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_123_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7895__A1 _2979_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6609_ _1745_ _1746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7589_ _2732_ _2736_ _2741_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_119_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5370__A2 _0497_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7647__A1 _2760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4881__A1 _3144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8503__C _3686_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4603__I net15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6689__A2 _1773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5361__A2 _0537_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7638__A1 _0940_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4872__A1 _4165_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6074__B1 _0052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6960_ _3926_ _2081_ _2083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5911_ _0703_ _1074_ _1075_ _1076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6891_ _2014_ _0014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8630_ _0104_ clknet_4_10_0_Clock C\[0\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5842_ _1004_ _1007_ _1008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6377__A1 _3999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8561_ _0006_ clknet_4_10_0_Clock A\[0\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5773_ _0937_ _0181_ _0920_ _0943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_72_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7512_ _2625_ _2626_ _2628_ _2662_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4724_ _3947_ _4045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_8492_ _3689_ _3690_ _0134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7877__A1 _2974_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7443_ _2469_ _2520_ _2590_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4655_ _3973_ _3976_ C\[3\]\[6\] _3977_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7374_ _2509_ _2514_ _2515_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4586_ _3901_ _3907_ _3908_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_11_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6325_ _1379_ _1473_ _1474_ _1475_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6256_ _1291_ _1332_ _1408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_118_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5207_ _2513_ _2599_ _0350_ _0388_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_88_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6852__A2 _1908_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6187_ _1227_ _1268_ _1343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4863__A1 _3971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8054__A1 _0633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5138_ _0319_ _0320_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6604__A2 _1740_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5069_ _0237_ _0245_ _0251_ _0252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_72_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6368__A1 _0062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6368__B2 _0063_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8109__A2 _3287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4423__I _2244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7580__A3 _1630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5591__A2 _0033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4394__A3 _3445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7868__A1 _0822_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6540__A1 _1619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5254__I B\[0\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7096__A2 _2170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5646__A3 _0451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6843__A2 _1968_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4854__A1 _3948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8045__A1 _1252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7020__A2 _1971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5031__A1 _0214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4333__I _2816_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8520__A2 _3687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4440_ B\[1\]\[1\] _3763_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4371_ _3218_ _3229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5164__I _0344_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6110_ _1225_ _1269_ _1270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_67_1366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7087__A2 _2188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7090_ _2176_ _2209_ _2210_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6041_ _1198_ _1203_ _1204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4845__A1 _4160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8036__A1 _0716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4508__I _3830_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6598__A1 _1732_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7992_ _0050_ _0013_ _3093_ _3162_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_81_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6943_ _3818_ _1907_ _2066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5270__A1 _0437_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6874_ _1998_ _1999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8613_ _0058_ clknet_4_1_0_Clock B\[3\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5825_ _4149_ _4189_ _0991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_22_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8544_ _3732_ _3734_ _3736_ _0146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5756_ _0024_ _0049_ _0926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4707_ _3841_ _3849_ _4028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8475_ _3673_ _3674_ _3675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5687_ _0858_ _0859_ _0860_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_124_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8511__A2 _3681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7426_ _2335_ _2485_ _2570_ _2571_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5325__A2 _0482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4638_ _3946_ _3960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_85_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7357_ _1247_ C\[1\]\[11\] _0476_ _2497_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4569_ _3890_ _3467_ _2764_ A\[3\]\[7\] _3891_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_104_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6308_ _1346_ _1387_ _1458_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7288_ _2349_ _2420_ _2421_ _2422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_81_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6239_ _1388_ _1391_ _1392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_77_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6825__A2 _1950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4836__A1 _4044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6589__A1 _1371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5958__B _0821_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6761__A1 _4076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4772__B1 _3893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8502__A2 _3676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6513__A1 _1604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6816__A2 _1922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4827__A1 _4127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8018__A1 _3186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5252__A1 _3892_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5004__A1 _0180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5610_ _0780_ _0782_ _0784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5555__A2 _0319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6590_ _1726_ _0000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6752__A1 _2449_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4998__I _4242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5541_ _0646_ _0718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8260_ _3394_ _3411_ _3453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_144_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6504__A1 _1590_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5472_ _0648_ _0649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7211_ _2334_ _2338_ _2339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_133_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4423_ _2244_ _3746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_126_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8191_ _0443_ _2045_ _3378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7142_ _2252_ _2263_ _2264_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4354_ _2503_ _3048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_141_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7073_ _2111_ _2193_ _2194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4285_ net1 _2319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4818__A1 _3111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8009__A1 _0319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6024_ _1175_ _1186_ _1187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__7480__A2 _0006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5491__A1 _0641_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4294__A2 _2405_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7232__A2 _2360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7975_ _0293_ _0298_ _0299_ _3146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6453__I _1597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6926_ _2046_ _2048_ _2049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_35_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8692__CLK clknet_4_5_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6857_ _3260_ _1848_ _1982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5808_ _0031_ _0057_ _4115_ _0974_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6788_ _3229_ _1811_ _1916_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8527_ _0131_ _3670_ _3721_ _0086_ _3722_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5739_ _0879_ _0880_ _0870_ _0911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_109_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7299__A2 _2257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8458_ _0937_ _3661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7409_ _3999_ _2404_ _2552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8389_ _3568_ _3573_ _3589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4809__A1 _4053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5482__A1 C\[2\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5482__B2 _3860_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4993__B1 _3391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5537__A2 _0711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7194__I _2234_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4611__I B\[1\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7143__B _2158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8565__CLK clknet_4_0_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5473__A1 _0386_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6017__A3 _4179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5225__A1 _0396_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7760_ _2914_ _2915_ _2916_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4972_ _0154_ _0156_ _0158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6711_ _1838_ _1841_ _1842_ _1843_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
X_7691_ _2806_ _2830_ _2843_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_1408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6642_ _1710_ _1777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5528__A2 _0393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6573_ _3531_ _1710_ _1711_ _1712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4521__I _3015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8312_ _3461_ _3477_ _3509_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_121_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5524_ _0699_ _0639_ _0700_ _0701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8243_ _3371_ _3433_ _3435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5455_ _0631_ _0632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7150__A1 _4090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4406_ _3551_ _3583_ _3593_ _3604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_8174_ _3299_ _3327_ _3360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5386_ _0511_ _0561_ _0562_ _0563_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5700__A2 _0462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4503__A3 _3825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7125_ _2147_ _2169_ _2247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4337_ _2856_ _2867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5352__I _0314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7056_ _2963_ _1863_ _2177_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_87_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5464__A1 _0629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6007_ _1026_ _1168_ _1169_ _1170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_67_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7205__A2 _1757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5301__B B\[0\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6559__A4 _2287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7756__A3 _2911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7958_ _0360_ _2077_ _3128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6909_ _1878_ _2031_ _2032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7889_ _3044_ _3043_ _3045_ _2970_ _3042_ _3052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_70_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4431__I _3753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8588__CLK clknet_4_2_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5207__A1 _2513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4606__I _3927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5758__A2 _0925_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6955__A1 _3832_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4430__A2 _3746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5930__A2 _1094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5143__B1 _0306_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5240_ _0419_ _0414_ _0420_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5171_ _0351_ _0352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_39_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput3 K[1] net3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_83_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7812_ _2904_ _2962_ _2969_ _2970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5749__A2 _3790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7743_ _2839_ _2892_ _2896_ _2898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4955_ _4265_ _4268_ _4269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8538__I2 _0105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7674_ _2825_ _2827_ _2828_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4886_ _3844_ _4202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6625_ _1745_ _1761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6556_ _1681_ _1683_ _1695_ _1697_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5507_ _0604_ _0621_ _0683_ _0684_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7123__A1 _2223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6487_ C\[2\]\[15\] _1630_ _1570_ _1631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8226_ _3359_ _3416_ _3417_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5438_ _3615_ _0363_ _0615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4488__A2 _3774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8157_ _3251_ _3252_ _3331_ _3341_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5369_ _0527_ _0545_ _0546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_82_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7108_ _2952_ _1927_ _2228_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7426__A2 _2485_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8088_ _3179_ _3263_ _3264_ _3265_ _3177_ _3266_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_82_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7039_ _4003_ _1791_ _2159_ _2160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_142_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5988__A2 _3872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6937__A1 _2042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7362__A1 _4069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5257__I _0435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7114__A1 _3861_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5125__B1 _0306_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7665__A2 _2776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4479__A2 net9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5720__I _0892_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8603__CLK clknet_4_0_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6928__A1 _3793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4740_ _4059_ _3769_ _4060_ _3770_ _4061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_124_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4671_ _3992_ _3993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7353__A1 _2430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6410_ _1554_ _1556_ _1557_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_70_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7390_ _2465_ _2530_ _2521_ _2531_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_70_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6341_ _1378_ _1382_ _1491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6272_ _1420_ _1421_ _1422_ _1423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_66_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7656__A2 _2777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8011_ _3181_ _3182_ _3183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5223_ _0356_ _0403_ _0404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7408__A2 _0005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5154_ _0335_ _0336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5085_ _0163_ _0164_ _0268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5987_ _2685_ _4135_ _1150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5198__A3 _0346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7592__A1 _2742_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4938_ _3944_ _4019_ _3913_ _4253_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_40_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7726_ _0775_ _1783_ _2882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7657_ _0752_ _1702_ _2810_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4869_ _4178_ _4184_ _4185_ _4186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_6608_ _3792_ _1744_ _1745_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7588_ _2740_ _0070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6539_ _1680_ _0124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5805__I _0220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7647__A2 _1762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8209_ _1178_ C\[0\]\[10\] _3398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8626__CLK clknet_4_2_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_7_0_Clock clknet_3_3_0_Clock clknet_4_7_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__4881__A2 _4196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6607__B1 _1743_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6636__I _1770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6083__A1 _1100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4872__A2 _4188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6074__A1 _3905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6074__B2 _3899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5910_ _0704_ _0705_ _1075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6890_ _2013_ _2014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5841_ _1002_ _1005_ _1006_ _1007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_22_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6377__A2 _0023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5772_ _0940_ _0941_ _0942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8560_ _0005_ clknet_4_10_0_Clock A\[0\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7511_ _2659_ _2660_ _2661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4723_ _3952_ _3953_ _3957_ _4044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_8491_ _0069_ _3687_ _3684_ _0065_ _3676_ _0067_ _3690_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_7442_ _2536_ _2587_ _2588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4654_ _3975_ _3976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7373_ _2510_ _2511_ _2512_ _2514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_4585_ _3902_ _3906_ _3907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8649__CLK clknet_4_11_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6324_ _1380_ _1381_ _1474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6255_ _1291_ _1332_ _1407_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_66_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5206_ _3531_ _2786_ _0330_ B\[0\]\[3\] _0387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_6186_ _1061_ _1224_ _1341_ _1342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4863__A2 C\[3\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8054__A2 _3104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5137_ _0318_ _0319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5360__I _0362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5068_ _0248_ _0249_ _0250_ _0251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA_input14_I Z[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5812__A1 _4127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6368__A2 _3900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7565__A1 _2646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5040__A2 _0222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7709_ _0761_ _1701_ _2863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8689_ _0135_ clknet_4_5_0_Clock net25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4394__A4 _3467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7868__A2 _2055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6540__A2 _1621_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4854__A2 _3936_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8045__A2 _1851_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6056__A1 _1057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5031__A2 _0208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4790__A1 _4025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7859__A2 _3018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4489__C _3701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4542__A1 _3860_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4370_ _3196_ _2405_ _3207_ _3218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6295__A1 _1428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6040_ _1199_ _1202_ _1203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I X[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8036__A2 _1715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6598__A2 _1734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7991_ _0052_ _1865_ _3003_ _3161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_54_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6942_ _3969_ _1726_ _2065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6873_ _1996_ _1997_ _3691_ _1998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_78_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8612_ _0057_ clknet_4_2_0_Clock B\[3\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5824_ _4165_ _4188_ _0990_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8543_ _0106_ _3714_ _3736_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5755_ _0903_ _0049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6770__A2 _1898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4706_ _2449_ _4026_ _4027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5686_ _0854_ _0855_ _0859_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8474_ _3664_ _3674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7425_ _0061_ _2014_ _2570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4637_ _3825_ _3951_ _3954_ _3958_ _3959_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_11_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4533__A1 _3854_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4568_ _2745_ _3890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7356_ _3998_ _2350_ _2496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6307_ _1457_ _0075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7287_ _2351_ _2353_ _2421_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4499_ _3821_ _3822_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6286__A1 _0456_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6238_ _1210_ _1389_ _1390_ _1391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6169_ _3961_ _1020_ _4096_ _1326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7786__A1 _2937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6589__A2 C\[1\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6210__A1 _1254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5564__A3 _0740_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6761__A2 _0001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4772__A1 B\[1\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4772__B2 _3783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5265__I _0325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7710__A1 _0335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4524__A1 _2971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4827__A2 _4144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4609__I _3916_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8018__A2 _3189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_4_0_Clock clknet_0_Clock clknet_3_4_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_48_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7777__A1 _2879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5252__A2 _0331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6752__A2 _1765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5540_ _4273_ _0716_ _0717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5471_ _0564_ _0565_ _3946_ _0648_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5175__I _3773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7701__A1 _2847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4422_ _3185_ net8 _3745_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4515__A1 _3037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7210_ _2335_ _2336_ _2337_ _2338_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_133_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8190_ _3374_ _3291_ _3376_ _3377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7141_ _2256_ _2262_ _2263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4353_ _2737_ _3037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__8501__I0 _0080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6268__A1 _3326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7072_ _2114_ _2192_ _2193_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_119_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4284_ B\[3\]\[2\] _2298_ _2308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_113_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4818__A2 _4135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6023_ _1177_ _1183_ _1185_ _1186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__8009__A2 _2045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5491__A2 _0645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7768__A1 _2870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4963__B _4276_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6734__I _1864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7974_ _3145_ _0114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6925_ _2031_ _2047_ _2048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_82_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6991__A2 _2093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6856_ _2492_ _1731_ A\[0\]\[5\] _1981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8193__A1 _0408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5807_ _4107_ _0031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5546__A3 _0722_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7940__A1 _0392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6787_ _1822_ _1828_ _1915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8601__D _0046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8526_ _3675_ _3668_ _3721_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5738_ _0902_ _0908_ _0909_ _0910_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4754__B2 _4044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8457_ _3660_ _0109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5669_ _3973_ C\[2\]\[1\] _0842_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_108_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7408_ _1530_ _0005_ _2551_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8388_ _3577_ _3579_ _3588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7339_ _2403_ _2408_ _2477_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6259__A1 _1167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4429__I B\[1\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5482__A2 _4242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7759__A1 _0838_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4993__A1 B\[1\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4993__B2 _3765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8184__A1 _3284_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5170__A1 _3456_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4339__I _2878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5473__A2 _4273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5225__A2 _0405_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4971_ _0154_ _0156_ _0157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_79_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6710_ _0513_ C\[1\]\[3\] _1842_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8175__A1 _3299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7690_ _2762_ _2840_ _2841_ _2842_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6641_ _3185_ _1733_ _1775_ _1776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7922__A1 _3960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4736__A1 _3955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6572_ A\[0\]\[0\] _1711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_125_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8311_ _3506_ _3507_ _3508_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5523_ _0637_ _0638_ _0700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5454_ _0630_ _0631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8242_ _3431_ _3432_ _3433_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4405_ _2674_ _3593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5385_ _0503_ _0560_ _0517_ _0562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_8173_ _3356_ _3357_ _3359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_99_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7124_ _2147_ _2169_ _2246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4336_ _2663_ _2856_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7055_ _2438_ _1927_ _2176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_86_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5464__A2 _0636_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6006_ _1028_ _1029_ _1031_ _1169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_95_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7957_ _0822_ _2185_ _3127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6908_ _3776_ _3004_ _1754_ _2031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_7888_ _3051_ _0128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6839_ _3004_ _1747_ _1965_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7913__A1 _3012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4712__I _3858_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4727__A1 _3932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8509_ _0097_ _0112_ _0082_ _0127_ _3704_ _3679_ _3706_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_104_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5543__I _0571_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5207__A2 _2599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6955__A2 _2077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4430__A3 _3747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7904__A1 _3792_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5930__A3 _0662_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5143__A1 net44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5143__B2 B\[2\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5170_ _3456_ _2816_ _0350_ _0351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8682__CLK clknet_4_11_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6643__A1 _3196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 K[2] net4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_65_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8396__A1 _3518_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7811_ _2906_ _2961_ _2969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_52_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6946__A2 _1993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5749__A3 _0920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7742_ _2842_ _2891_ _2896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4957__A1 _3814_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4954_ _4266_ _4267_ _4268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8538__I3 _0090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7673_ _0035_ _1716_ _2824_ _1534_ _2827_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_71_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4885_ _3056_ _3089_ _3794_ _4200_ _4201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_123_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6624_ _3904_ _1740_ _1749_ _1759_ _1760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_53_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6555_ _1681_ _1683_ _1695_ _1696_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_69_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5506_ _0606_ _0620_ _0683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7659__B1 _1747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6486_ _1534_ _1630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5134__A1 _0310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8225_ _3362_ _3415_ _3416_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_106_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5437_ _0612_ _0542_ _0613_ _0614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6882__A1 _1939_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5368_ _0528_ _0544_ _0545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8156_ _3251_ _3252_ _3331_ _3340_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7107_ _3015_ _1863_ _2227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4319_ _2545_ _2642_ _2674_ _2685_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_5299_ _4130_ _0472_ _0474_ _0476_ _0477_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8087_ _3179_ _3193_ _3265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7426__A3 _2570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6634__A1 _1768_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7038_ _4089_ C\[1\]\[7\] _2159_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6194__I _0687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8555__CLK clknet_4_2_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4442__I _3755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_4_3_0_Clock clknet_3_1_0_Clock clknet_4_3_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__7362__A2 _1529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7114__A2 _1808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5125__A1 _3271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5125__B2 B\[2\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5676__A2 _0847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7702__B _2829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6928__A2 _3861_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4352__I _3015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4670_ _3991_ _3992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6340_ _1475_ _1489_ _1490_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8302__A1 _0053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6271_ _3883_ _3899_ _1422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5183__I _0363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6864__A1 _1984_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5222_ _0391_ _0403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8010_ _0529_ _1928_ _3182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8494__I _3692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5153_ _3778_ _0335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_111_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5084_ _0264_ _0265_ _0266_ _0267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4627__B1 _3271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6631__A4 _1765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8578__CLK clknet_4_1_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6919__A2 _1968_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7041__A1 _1018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5986_ _1147_ _1148_ _1149_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7592__A2 _2743_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7725_ _0488_ _2771_ _2881_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4937_ _4236_ _4250_ _4251_ _4252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7656_ _2770_ _2777_ _2809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4868_ _3793_ _3937_ _3980_ _4185_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_36_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5355__A1 _0440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6607_ _3797_ _1742_ _1743_ A\[1\]\[1\] _1744_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_7587_ _0950_ _0951_ _2740_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4799_ _4116_ _4117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6538_ _1670_ _1679_ _1680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_14_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5107__A1 _0285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6469_ _1613_ _1548_ _1614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7647__A3 _1814_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5658__A2 _0830_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8208_ _3395_ _3317_ _3396_ _3397_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4866__B1 _4180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8139_ _3220_ _3223_ _3322_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6607__A1 _3797_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6607__B2 A\[1\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6083__A2 _1102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4437__I _3759_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7280__A1 _2411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7032__A1 _4150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5594__A1 _2889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8532__A1 _3692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5897__A2 _1060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4900__I _4214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5731__I _0493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6074__A2 _0053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5282__B1 _0306_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6562__I _1701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5840_ _0800_ _3873_ _1006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5585__A1 _3876_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5771_ _0928_ _0929_ _0921_ _0941_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_99_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7510_ _4035_ _2390_ _2616_ _2660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4722_ _3988_ _4018_ _4042_ _4043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8490_ _0071_ _3669_ _3689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7441_ _2539_ _2586_ _2587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4653_ _3974_ _3975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7372_ _1538_ _0005_ _2512_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4584_ _3904_ _3905_ _3906_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6323_ _1380_ _1381_ _1473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6837__A1 _4007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6254_ _1147_ _1287_ _1406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5205_ _3956_ _0386_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6185_ _1216_ _1340_ _1341_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5136_ _0317_ _0318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7262__A1 _2346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5067_ _0025_ _4117_ _4263_ _0205_ _0250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_85_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5812__A2 _4144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8604__D _0049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5969_ _0994_ _0995_ _1010_ _1133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7708_ _0751_ _1746_ _2862_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8688_ _0134_ clknet_4_5_0_Clock net24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7317__A2 _2377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5328__A1 _2755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7639_ _0941_ _2790_ _2791_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_119_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6056__A2 _1079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7253__A1 _2309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6382__I _1529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8505__A1 _3702_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5319__A1 _4072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_0_0_Clock clknet_0_Clock clknet_3_0_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_89_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4630__I _3761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4542__A2 _3864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8036__A3 _3112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7990_ _3000_ _3082_ _3159_ _3098_ _3087_ _3160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_93_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5255__B1 _0432_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7795__A2 _4239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6941_ _1979_ _2061_ _2062_ _2002_ _2043_ _2063_ _2064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai33_1
XFILLER_82_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6872_ _3802_ _1710_ _1997_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8611_ _0056_ clknet_4_1_0_Clock B\[3\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5823_ _4165_ _4188_ _0989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_50_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8542_ _3693_ _3733_ _3708_ _3734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5754_ _0924_ _0925_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8616__CLK clknet_4_1_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4705_ _3304_ _4026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8473_ net14 _3673_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4781__A2 _4100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5685_ _0857_ _0858_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4540__I _3862_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7424_ _2548_ _2568_ _2569_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4636_ _3955_ _3956_ _3957_ _3958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_50_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4533__A2 _3467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7355_ _2439_ _2442_ _2494_ _2495_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4567_ _3888_ _3889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6306_ _1405_ _1456_ _1457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_85_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7286_ _2351_ _2353_ _2420_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4498_ _2867_ _3821_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6286__A2 C\[3\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6237_ _1213_ _1270_ _1390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6168_ _1323_ _1324_ _1325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7235__A1 _3957_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5119_ _4261_ _0301_ _0302_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_79_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6099_ _1245_ _1258_ _1259_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_58_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6589__A3 _1723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6930__I _4214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6210__A2 _1255_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8499__B1 _3697_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4772__A2 _3780_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4450__I _3772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7710__A2 _0896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4524__A2 _3846_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5721__A1 _0336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7474__A1 _1533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5788__A1 _0914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4625__I _3946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4460__A1 _2352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8639__CLK clknet_4_2_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7157__B _3991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5960__A1 _1121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5456__I _0568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5470_ _0646_ _0647_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4421_ _3735_ _3744_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4515__A2 _3048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7140_ _2260_ _2261_ _2262_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4352_ _3015_ _3026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6268__A2 _1419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7465__A1 _1419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7071_ _2130_ _2132_ _2191_ _2192_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_4283_ _2233_ _2254_ _2276_ _2287_ _2298_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_80_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6022_ _1184_ _4080_ _4096_ _1185_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_98_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7768__A2 _2877_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7973_ _3052_ _3143_ _3145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_54_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6924_ _3792_ _2941_ _1807_ _2047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_81_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6855_ _1971_ _1980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_126_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8193__A2 _1929_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5806_ _4107_ _0057_ _4115_ _0973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_11_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6786_ _0202_ _1763_ _0011_ _1914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_91_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7940__A2 _2250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8525_ _3719_ _0101_ _3720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5951__A1 _1051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5737_ _0906_ _0907_ _0909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4754__A2 _4068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8456_ _3649_ _3655_ _3659_ _3660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_108_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5668_ _0776_ _0840_ _0841_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7407_ _2436_ _2499_ _2549_ _2550_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5703__A1 _0200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4506__A2 net10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4619_ _3939_ _3940_ _3941_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8387_ _3587_ _0106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5599_ _0763_ _0771_ _0772_ _0773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7338_ _2417_ _2446_ _2475_ _2476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7456__A1 _2485_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7269_ _4133_ _1864_ _2401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7208__A1 _4133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7759__A2 _2120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4445__I A\[2\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4993__A2 _3764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6195__A1 _0030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5942__A1 _0422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5170__A2 _2816_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7998__A2 _3109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5473__A3 _0647_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4970_ _0155_ _4210_ _0156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_45_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8702__D _0148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6640_ A\[0\]\[1\] _1775_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_75_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7922__A2 _0325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6571_ _1709_ _1710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4736__A2 _4009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8310_ _3503_ _3505_ _3507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5522_ _0637_ _0638_ _0699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8241_ _3366_ _3385_ _3432_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5453_ _0564_ _0565_ _0630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7150__A3 _2156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4404_ _2794_ _2836_ _3572_ _3583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_8172_ _0897_ _2390_ _3285_ _3284_ _3267_ _3357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_99_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5384_ _0560_ _0517_ _0503_ _0561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7123_ _2223_ _2243_ _2245_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4335_ _2794_ _2826_ _2836_ _2845_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7989__A2 _3098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7054_ _3991_ _2993_ _1807_ _2175_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_87_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6005_ _1028_ _1029_ _1031_ _1168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_132_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4672__A1 _3993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7956_ _3123_ _3124_ _3125_ _3126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6907_ _1965_ _1967_ _2030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7887_ _3050_ _0961_ _3051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_126_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8612__D _0057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6838_ _1961_ _1963_ _1964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7913__A2 _3038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4727__A2 _4044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6769_ _3819_ _1733_ _1898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8508_ _3705_ _0137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8439_ _3627_ _3630_ _3642_ _3643_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_137_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6101__A1 _1105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4663__A1 _3979_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4415__A1 _2481_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4966__A2 _0151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4903__I _4071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7904__A2 _0317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5391__A2 _0505_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7668__A1 _0435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5143__A2 _0304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6340__A1 _1475_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8093__A1 _3198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6643__A2 _1777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7840__A1 _0344_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput5 X[0] net5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8396__A2 _0007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7810_ _2968_ _0127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4406__A1 _3551_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7741_ _2895_ _0126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4953_ _0028_ _3889_ _4267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4957__A2 _4007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8148__A2 _3331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7672_ _0035_ _1716_ _2824_ _2825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_75_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4884_ _2941_ _4200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6623_ _1758_ _1759_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6554_ _1686_ _1691_ _1694_ _1695_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__5382__A2 _0558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5505_ _0589_ _0593_ _0682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7659__A1 _0752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7659__B2 _0896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6485_ C\[2\]\[15\] _1628_ _1629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_134_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8224_ _3386_ _3414_ _3415_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_10_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5436_ _4173_ _4026_ _0364_ _0355_ _0613_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_133_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5134__A2 _0315_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6331__A1 _1374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8155_ _3052_ _3141_ _3244_ _3140_ _3339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_5367_ _0532_ _0536_ _0543_ _0544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_114_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4893__A1 _0028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7106_ _4112_ _2012_ _2226_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4318_ _2663_ _2674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_8086_ _3184_ _3192_ _3264_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_101_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5298_ _3974_ _0476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7037_ _2084_ _2088_ _2157_ _2158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6634__A2 _1702_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8607__D _0052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4645__A1 _3413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6398__A1 _1429_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7939_ _3105_ _3106_ _3107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7362__A3 _0004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6570__A1 net3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5125__A2 _0304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5676__A3 _0848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5503__B _0670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7822__A1 _1753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4636__A1 _3955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6389__A1 _0337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6928__A3 _2050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7050__A2 _2057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4633__I _3709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7889__B2 _3042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8302__A2 _2203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6270_ _0062_ _3905_ _1421_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5221_ _4213_ _0401_ _0402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6864__A2 _1988_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5152_ _0333_ _0334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5083_ _0238_ _0241_ _0266_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4627__A1 B\[1\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4627__B2 _3783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5985_ _4195_ _3897_ _3625_ _4202_ _1148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7724_ _0035_ _1716_ _2824_ _2880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_75_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4936_ _4248_ _4249_ _4251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7655_ _2807_ _2778_ _2808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4867_ _4181_ _4183_ _4184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6606_ _3358_ _3779_ _2373_ _2567_ _1743_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7586_ _2739_ _0064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4798_ _3903_ _4116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6537_ _1639_ _1675_ _1678_ _1679_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_105_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6468_ _1511_ _1613_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8207_ _3312_ _3314_ _3396_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5419_ _0527_ _0545_ _0596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6399_ _1544_ _1545_ _1546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4866__A1 _3777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4866__B2 _4087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8138_ _3221_ _3222_ _3321_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6607__A2 _1742_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8069_ _3244_ _3246_ _3247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_130_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4618__A1 C\[3\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6083__A3 _1103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7280__A2 _2412_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7032__A2 _2152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4453__I _3775_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8672__CLK clknet_4_4_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6791__A1 _3888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5594__A2 _0363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5284__I _0461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4857__A1 _0043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4628__I _3949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7271__A2 _2402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5282__A1 _0430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5282__B2 _0459_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5770_ _0937_ _0181_ _0920_ _0939_ _0940_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_61_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5585__A2 _0315_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6782__A1 _1893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4721_ _3945_ _3987_ _4042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7440_ _2542_ _2585_ _2586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4652_ _2652_ _3974_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7371_ _2087_ _0005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4583_ _3636_ _3905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6322_ _1351_ _1471_ _1472_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_115_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6253_ _1400_ _1404_ _1405_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6837__A2 _1962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4848__A1 _4095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5204_ _0374_ _0378_ _0384_ _3997_ _0385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6184_ _1223_ _1340_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5135_ _3819_ net45 _0312_ B\[2\]\[4\] _0317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_135_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5066_ _0027_ _0056_ _0220_ _0026_ _0249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5273__A1 _0340_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8695__CLK clknet_4_7_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8211__A1 _0630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5025__A1 _0025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5968_ _0998_ _1009_ _1132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4919_ _4233_ _4234_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7707_ _2859_ _2860_ _2825_ _2827_ _2861_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_8687_ _0133_ clknet_4_5_0_Clock net16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5899_ _1055_ _1063_ _1064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_138_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8620__D _0069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7638_ _0940_ _0953_ _2790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5328__A2 _3562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5879__A3 _1044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7569_ _1688_ C\[1\]\[16\] _2723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8278__A1 _3465_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7789__B1 _1972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8202__A1 _3305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5279__I _0456_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5319__A2 _0393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7713__B1 _0002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8269__A1 _3462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8568__CLK clknet_4_3_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5255__A1 _0430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6940_ _1974_ _1976_ _2063_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_81_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6871_ _2330_ _1707_ _1995_ _1996_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5007__A1 _4270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5822_ _0973_ _0987_ _0988_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8610_ _0055_ clknet_4_11_0_Clock B\[2\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5558__A2 _0734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8541_ _0121_ _0076_ _3695_ _3733_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5753_ _0922_ _0923_ _0924_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4704_ _3996_ _4023_ _4024_ _4025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8472_ _1696_ _1697_ _3670_ _3671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5684_ _0835_ _0836_ _0857_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_120_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7423_ _2558_ _2566_ _2568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4635_ _3934_ _3957_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_141_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7354_ _2367_ _2437_ _2494_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_116_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4566_ _3499_ _3888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4533__A3 _2764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6305_ _1451_ _1455_ _1456_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_131_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7285_ _2355_ _2371_ _2418_ _2419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4497_ B\[1\]\[4\] _3781_ _3819_ _3784_ _3820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_143_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6236_ _1213_ _1270_ _1389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6167_ _3961_ _4079_ _4093_ _1322_ _4088_ _1324_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
XTAP_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5118_ _0178_ _0300_ _0301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6098_ _1246_ _1251_ _1257_ _1258_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_3517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6589__A4 _1726_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8615__D _0060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5049_ _0191_ _0198_ _0232_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_45_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6994__A1 _0202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5549__A2 _0618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6746__A1 _1832_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8499__A1 _0102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8499__B2 _0072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7710__A3 _2237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5721__A2 _0334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7474__A2 _1983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5485__A1 _3972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5237__A1 _4073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4996__B1 _4150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8187__B1 _1810_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4460__A2 _3748_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6737__A1 _0057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5960__A2 _1124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4420_ _2737_ _3727_ _2373_ _2503_ _3735_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__5712__A2 _0884_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4351_ _3004_ _3015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5472__I _0648_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7070_ _2135_ _2170_ _2190_ _2191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__7465__A2 _2579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4282_ net4 _2287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_113_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6021_ _3992_ _1184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6425__B1 _1094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5779__A2 _0947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7972_ _3140_ _3142_ _3143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6923_ _4112_ _2045_ _2046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4451__A2 _3767_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6854_ _1901_ _1977_ _1978_ _1979_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_1440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5805_ _0220_ _0057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6785_ _1812_ _0011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4551__I _3873_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8524_ _3683_ _3719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5736_ _0906_ _0907_ _0908_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_109_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5667_ _0839_ _0840_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7153__A1 _3982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8455_ _3630_ _3656_ _3657_ _3658_ _3659_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_50_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7406_ _2500_ _2505_ _2549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4618_ C\[3\]\[5\] _3928_ _3940_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8386_ _3584_ _3586_ _3587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5703__A2 _0838_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5598_ _0767_ _0770_ _0772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7337_ _2419_ _2445_ _2475_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4549_ _3867_ _3872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7268_ _2348_ _2398_ _2399_ _2400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6219_ _1247_ _1374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7199_ _2256_ _2262_ _2326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_131_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7208__A2 _1809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8405__A1 _3553_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5219__A1 _0379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4690__A2 _4009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5331__B _3990_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6719__A1 _1847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6195__A2 _0054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4461__I _3783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5942__A2 _0720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7144__A1 _2158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5155__B1 net44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7695__A2 _2777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5458__A1 _3965_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8606__CLK clknet_4_1_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6958__A1 _1178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7922__A3 _2050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6570_ net3 net2 net4 _1709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__5933__A2 _0722_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4736__A3 _4056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5521_ _0641_ _0696_ _0697_ _0698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8240_ _3368_ _3384_ _3431_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5452_ _0626_ _0627_ _0628_ _0629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5697__A1 _0753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4403_ _3562_ _3572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_8171_ _3278_ _3295_ _3355_ _3356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5383_ _0516_ _0560_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_126_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7122_ _2225_ _2242_ _2243_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4334_ _2621_ _2836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_99_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7053_ _1984_ _2067_ _2174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6004_ _1165_ _1166_ _1167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4672__A2 _3786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7955_ _3013_ _3014_ _3125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6906_ _1960_ _1969_ _2029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7886_ _0918_ _0960_ _3050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6837_ _4007_ _1962_ _1963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7374__A1 _2509_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4281__I _2265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6768_ _3542_ _1777_ A\[0\]\[4\] _1897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8507_ _0096_ _0111_ _0081_ _0126_ _3704_ _3679_ _3705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5719_ _0888_ _0891_ _0892_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_52_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6699_ _1795_ _1793_ _1831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8438_ _3631_ _3641_ _3642_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_136_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8369_ _1094_ _0055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6001__I _1163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8629__CLK clknet_4_8_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4360__A1 _3056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6101__A2 _1106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5860__A1 _4183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4663__A2 _3981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4456__I _3727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5612__A1 _0022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4415__A2 net15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8157__A3 _3331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7904__A3 _3002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7117__A1 _2236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7668__A2 _0003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8547__B _3708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6846__I _1971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5750__I _0774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7840__A2 _1863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput6 X[1] net6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6800__B1 _1698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7740_ _0956_ _0957_ _2895_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_64_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4952_ _4263_ _4264_ _4266_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_51_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4883_ _2460_ _4198_ _4199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5197__I _0377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7356__A1 _3998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7671_ _1479_ C\[0\]\[3\] _2824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6622_ _1757_ _1758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6553_ _1655_ _1662_ _1692_ _1653_ _1693_ _1694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_5504_ _0599_ _0671_ _0680_ _0681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4590__A1 _3682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6484_ _0947_ _1628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7659__A2 _1703_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8223_ _3388_ _3412_ _3414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_69_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5435_ _4026_ _0364_ _0355_ _0422_ _0612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_105_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6331__A2 C\[2\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8154_ _3338_ _0116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5366_ _0538_ _0540_ _0542_ _0543_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_142_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6882__A3 _2006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4893__A2 _3240_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7105_ _2136_ _2143_ _2224_ _2225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4317_ _2319_ _2652_ _2663_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_113_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8085_ _3184_ _3192_ _3263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5297_ _3304_ _0472_ _0474_ _0475_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_114_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6095__A1 _3831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7036_ _1372_ C\[1\]\[6\] _2156_ _1826_ _2157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_45_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4645__A2 net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7595__A1 _2733_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8623__D _0111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7938_ _0481_ _1841_ _1903_ _0382_ _3106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7869_ _0924_ _2257_ _3033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7347__A1 _3877_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7362__A4 _2501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6570__A2 net2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7822__A2 _0317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5833__A1 _2460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4636__A2 _3956_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6389__A2 _1533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5061__A2 _0243_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6010__A1 _0021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8121__I _2077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7510__A1 _4035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5220_ _0400_ _0401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5151_ _3892_ _3391_ _0331_ _0332_ B\[0\]\[0\] _0333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_97_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5480__I _0656_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7813__A2 _2918_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5082_ _0238_ _0241_ _0265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5824__A1 _4165_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4627__A2 _3780_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5984_ _1000_ _1146_ _1147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7723_ _2870_ _2877_ _2879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7329__A1 _2385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4935_ _4248_ _4249_ _4250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7654_ _2770_ _2777_ _2807_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4866_ _3777_ _3823_ _4182_ _4180_ _4087_ _4183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_6605_ _3746_ _3748_ _2394_ _1742_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_123_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4797_ _3846_ _4028_ _4114_ _4115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7585_ _0209_ _0224_ _2739_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4563__A1 _3882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6536_ _1676_ _1637_ _1677_ _1678_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6467_ _1591_ _1611_ _1612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_133_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8206_ _0632_ _1975_ _3313_ _3395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4315__A1 _2578_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5418_ _0528_ _0544_ _0595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6398_ _1429_ _1444_ _1545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4866__A2 _3823_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6486__I _1534_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8618__D _0063_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5349_ _0418_ _0425_ _0526_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8137_ _3301_ _3319_ _3320_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_87_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8068_ _3142_ _3245_ _3246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4618__A2 _3928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7019_ _3816_ _2139_ _2140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7568__A1 _2659_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5579__B1 _3271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6791__A2 _1865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4306__A1 _2492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4857__A2 _4173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5806__A1 _4107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5282__A2 _0304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4644__I B\[1\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6231__A1 _1365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6782__A2 _1910_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4720_ _3880_ _4040_ _4041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4651_ _3972_ _3973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7731__A1 _2861_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4545__A1 _3867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4582_ _3903_ _3904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7370_ _1295_ _1949_ _2511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6321_ _0327_ _1357_ _1358_ _1470_ _1471_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__8531__I0 _0118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6252_ _1194_ _1197_ _1402_ _1403_ _1404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_115_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5203_ _0383_ _0384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4848__A2 _4097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4819__I _4135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6183_ _1339_ _0074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5134_ _0310_ _0315_ _0316_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5065_ _0247_ _0248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4554__I _3864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8211__A2 _2275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5025__A2 _0202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5967_ _0988_ _1129_ _1130_ _1131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_52_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7706_ _2819_ _2823_ _2860_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4918_ _4212_ _4230_ _4233_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8686_ _0079_ clknet_4_13_0_Clock C\[3\]\[16\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5898_ _1061_ _1062_ _1063_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7637_ _2789_ _0072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5328__A3 _0380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4849_ _3970_ _3984_ _4166_ _4098_ _4083_ _4167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_53_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7568_ _2659_ _2711_ _2709_ _2722_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6519_ _1515_ _1661_ _1662_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_88_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8522__I0 _0085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7499_ _2648_ _0091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6289__A1 _1438_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6461__A1 _1604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4472__B1 _2897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6213__A1 _1246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7961__A1 _3126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4775__A1 _4086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5295__I _4089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6516__A2 _0947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7713__A1 _0899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7713__B2 _0925_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4527__A1 _3848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4527__B2 _3849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8269__A2 _0003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4639__I _3960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6870_ A\[0\]\[4\] _1995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5007__A2 _4271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5821_ _0985_ _0986_ _0987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_62_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8540_ _0091_ _3676_ _3732_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4766__A1 _3983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5752_ _0359_ _0923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4703_ _4000_ _4005_ _4017_ _4024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8471_ _3668_ _3670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6507__A2 _1615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5683_ _0854_ _0855_ _0856_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7422_ _2559_ _2565_ _2566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4634_ _3920_ _3956_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7180__A2 _2288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5191__A1 _0366_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4565_ _3837_ _3880_ _3881_ _3885_ _3886_ _3887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_7353_ _2430_ _2444_ _2491_ _2493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6304_ _1453_ _1454_ _1455_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_144_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4496_ _2982_ _3819_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7284_ _2358_ _2370_ _2418_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4549__I _3867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6235_ _1342_ _1346_ _1387_ _1388_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_131_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8662__CLK clknet_4_14_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5494__A2 _0670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6691__A1 _4200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6166_ _1184_ _4079_ _4176_ _1322_ _1323_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_1
XTAP_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5117_ _0176_ _0177_ _0293_ _0298_ _0299_ _0300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_2
XTAP_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8432__A2 _1628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6097_ _1253_ _1256_ _1257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_100_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5246__A2 _0418_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5048_ _0218_ _0230_ _0231_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_22_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input12_I X[7] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6994__A2 _0013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7943__A1 _3423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6746__A2 _1854_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6999_ _1949_ _2120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8631__D _0105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8499__A2 _3666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8669_ _0124_ clknet_4_15_0_Clock C\[2\]\[16\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5485__A2 C\[2\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6682__A1 _4116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4693__B1 _3967_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4996__A1 _3979_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4996__B2 _0181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8187__A1 _1099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8187__B2 _0444_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4460__A3 _3782_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6737__A2 _0008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6849__I _1839_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8685__CLK clknet_4_13_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4350_ _2993_ _3004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4920__A1 _4224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8111__A1 _0409_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4281_ _2265_ _2276_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_119_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6020_ _1180_ _1182_ _1183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input4_I K[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6425__A1 C\[2\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6425__B2 _3898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7971_ _3141_ _3142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6976__A2 _3709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6922_ _1862_ _2045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4451__A3 _3773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6853_ _1895_ _1906_ _1908_ _1978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_63_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7925__A1 _0314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5804_ _3911_ _4193_ _0971_ _0972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__4739__A1 _3423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6784_ _1887_ _1889_ _1912_ _1913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_8523_ _3717_ _0141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5735_ _0848_ _0876_ _0877_ _0907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_50_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8454_ _3631_ _3641_ _3658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5666_ _0203_ _0838_ _0775_ _0774_ _0839_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7405_ _2546_ _2547_ _2548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4617_ _3932_ _3935_ _3938_ _3939_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_135_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8385_ _3539_ _3541_ _3585_ _3586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5597_ _0767_ _0770_ _0771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_89_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4911__A1 _4224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7336_ _2411_ _2473_ _2474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_85_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4548_ _3870_ _3871_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8102__A1 _3201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4279__I _2244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7267_ _2270_ _2354_ _2399_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4479_ _2233_ net9 _3802_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_131_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6218_ _1372_ C\[2\]\[12\] _0469_ _1373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_58_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7198_ _2322_ _2324_ _2325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8626__D _0114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6149_ _0021_ _3999_ _1174_ _1308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5219__A2 _0381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4690__A3 _4010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4978__A1 _4238_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8558__CLK clknet_4_8_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6719__A2 _1850_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8341__A1 _3427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5155__A1 A\[2\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5155__B2 _4077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7695__A3 _2813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4902__A1 _3774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5458__A2 _4213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7852__B1 _2871_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6958__A2 C\[1\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4969__A1 _4227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5748__I _0334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7907__A1 _0903_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4652__I _2652_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_0_0_Clock_I clknet_3_0_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5520_ _0645_ _0667_ _0697_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5451_ _0554_ _0555_ _0628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4402_ _2330_ net11 _3562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_4
X_8170_ _3281_ _3294_ _3355_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5382_ _0552_ _0558_ _0559_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_126_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7121_ _2230_ _2234_ _2241_ _2242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_86_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4333_ _2816_ _2826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_99_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7052_ _2049_ _2171_ _2172_ _2173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6003_ _1022_ _1023_ _1166_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8399__A1 _1673_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8700__CLK clknet_4_13_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7954_ _0389_ _1962_ _3124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7359__B _2498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6905_ _2026_ _2027_ _2028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_82_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7885_ _3049_ _0083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6836_ _1902_ _1962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6767_ _3931_ _1725_ _1896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8506_ _3674_ _3704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_13_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5718_ _0889_ _0890_ _0861_ _0891_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_137_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8323__A1 _0457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6698_ _1829_ _1830_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8437_ _3591_ _3640_ _3641_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5649_ _0347_ _0351_ _0822_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8368_ _3497_ _3502_ _3568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7319_ _2452_ _2455_ _2456_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4360__A2 _3089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8299_ _3494_ _3490_ _3495_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7062__A1 _3960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5612__A2 _0436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5915__A3 _1079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7117__A2 _2179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6876__A1 _1905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6628__A1 _0208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4647__I _3968_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput7 X[2] net7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7053__A1 _1984_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6862__I _1986_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5603__A2 _0493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6800__A1 _1926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6800__B2 _3829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4951_ _4263_ _4264_ _4265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7670_ _0403_ _0035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4882_ _3848_ _4198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8553__A1 _3645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7356__A2 _2350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6621_ _1756_ _1757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6552_ _1651_ _1663_ _1693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_119_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7108__A2 _1927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8305__A1 _3498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5503_ _0600_ _0679_ _0670_ _0680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6483_ _1564_ _1579_ _1627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6867__A1 _4087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8222_ _3390_ _3394_ _3411_ _3412_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_5434_ _0608_ _0610_ _0611_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_133_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6331__A3 B\[2\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8153_ _3332_ _3336_ _3338_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_86_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5365_ _0541_ _0423_ _0542_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7104_ _2137_ _2142_ _2224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4316_ net15 _2652_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8084_ _3161_ _3162_ _3165_ _3262_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5296_ _0473_ C\[2\]\[5\] _0474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6095__A2 _0569_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7035_ _2155_ _2156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7044__A1 _1838_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7937_ _0382_ _0509_ _3104_ _2275_ _3105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_93_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4292__I _2383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7868_ _0822_ _2055_ _3032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7347__A2 _2120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6819_ _1880_ _1886_ _1945_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5358__A1 _3806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7799_ _2935_ _2958_ _2959_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6570__A3 net4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7283__A1 _2397_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4467__I _3789_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7822__A3 _1755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5833__A2 _3897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4636__A3 _3957_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5349__A1 _0418_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6010__A2 _3998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7510__A2 _2390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5521__A1 _0641_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5150_ _3982_ _3892_ _0331_ _0332_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_69_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7274__A1 _2053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5081_ _0244_ _0264_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5824__A2 _4188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7026__A1 _2137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7026__B2 _2080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5983_ _3844_ _0574_ _1146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7722_ _2875_ _2876_ _2877_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_80_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4934_ _3930_ _3941_ _3914_ _4249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__8619__CLK clknet_4_1_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8526__A1 _3675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7653_ _0897_ _1704_ _2803_ _2804_ _2806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4865_ _4092_ _4182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4840__I _4066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6604_ _0211_ _1740_ _1741_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7584_ _2738_ _0068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4796_ _0058_ _0029_ _4029_ _4114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_105_1440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6535_ _1632_ _1634_ _1677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5760__A1 _0928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4563__A2 _0061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6466_ _1608_ _1610_ _1611_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_49_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8205_ _3308_ _3392_ _3393_ _3394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5417_ _0589_ _0593_ _0594_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4315__A2 _2599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6397_ _1433_ _1443_ _1544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8136_ _3308_ _3311_ _3318_ _3319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_87_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4866__A3 _4182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5348_ _0418_ _0425_ _0525_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8067_ _3052_ _3140_ _3245_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5279_ _0456_ _0457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7018_ _2054_ _2139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7017__A1 _4135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5579__A1 A\[2\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5579__B2 _4077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8517__A1 _3692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4750__I _3751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5067__B _4263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6677__I _1809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4306__A2 _2513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5806__A2 _0057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5990__A1 _3862_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4660__I _3890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4650_ _3971_ _3972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput10 X[5] net10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5742__A1 _0895_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4545__A2 _3122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4581_ _3229_ _3903_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6320_ _1357_ _1358_ _1469_ _1470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8531__I1 _0073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6251_ _1280_ _1401_ _1335_ _1403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5202_ _0382_ _0383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_103_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6182_ _1336_ _1338_ _1339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_135_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5133_ _0314_ _0315_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5064_ _0205_ _0246_ _0212_ _0247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_69_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4481__A1 _3802_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6222__A2 _1376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5966_ _0993_ _1044_ _1130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_53_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7705_ _2819_ _2823_ _2859_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_80_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4917_ _4212_ _4230_ _4231_ _4232_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8685_ _0078_ clknet_4_13_0_Clock C\[3\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5981__A1 _4215_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5897_ _1059_ _1060_ _1062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8591__CLK clknet_4_9_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7636_ _0218_ _2788_ _2789_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_107_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4848_ _4095_ _4097_ _4166_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_119_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5733__A1 _0847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7567_ _2682_ _2719_ _2720_ _2715_ _2721_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_1210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4779_ _4083_ _4098_ _4099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_101_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6518_ _1656_ _1660_ _1661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_4_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7498_ _2640_ _2644_ _2647_ _2648_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_107_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8522__I1 _0100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8629__D _0103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6449_ _1592_ _1593_ _1594_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_134_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8119_ _3225_ _3232_ _3300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_76_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7789__A2 _1771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4745__I _3821_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4472__B2 _3788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5972__A1 _0060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5576__I _0751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4480__I A\[2\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7713__A2 _0001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4527__A2 _3026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7229__A1 _2269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6204__A2 _1358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6870__I A\[0\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7401__A1 _2490_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5007__A3 _4274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5820_ _0978_ _0979_ _0984_ _0986_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_50_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5751_ _0358_ _0922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_97_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5963__A1 _0973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4766__A2 C\[3\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4390__I _3423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4702_ _4000_ _4005_ _4017_ _4023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8470_ _3668_ _3669_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5682_ _0790_ _0806_ _0855_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_124_1156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7421_ _2560_ _2564_ _2565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5715__A1 _0867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4633_ _3709_ _3955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7352_ _2433_ _2443_ _2491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5191__A2 _0370_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4564_ _3837_ _3852_ _3879_ _3886_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_50_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6303_ _1282_ _1334_ _1454_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7283_ _2397_ _2415_ _2417_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_85_1449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4495_ _3817_ _3818_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6234_ _1354_ _1386_ _1387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6140__A1 _3883_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6691__A2 _1823_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6165_ _0473_ C\[3\]\[11\] _1322_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5116_ _0296_ _0297_ _0299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_85_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6096_ _1254_ _1255_ _1256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_131_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5246__A3 _0425_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5047_ _0219_ _0229_ _0230_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5651__B1 _0823_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6998_ _2031_ _2047_ _2119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5949_ _1065_ _1069_ _1113_ _1114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_40_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8668_ _0123_ clknet_4_15_0_Clock C\[2\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7619_ _1713_ _2771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8599_ _0044_ clknet_4_3_0_Clock B\[1\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7459__A1 _2603_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6682__A2 _0009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4693__B2 _3770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5237__A3 _0414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4996__A2 _3799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8187__A2 _1765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6690__I _1700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7719__C _4066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7934__A2 _2955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5945__A1 _1098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_3_0_0_Clock_I clknet_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_118_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4920__A2 _4225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8111__A2 _1864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4280_ net2 _2265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_49_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7870__A1 _0435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7622__A1 _2773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6425__A2 _0185_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7970_ _3054_ _3057_ _3139_ _3141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6976__A3 _1743_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6921_ _1961_ _1963_ _2044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6852_ _1906_ _1908_ _1895_ _1977_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5803_ _4105_ _4192_ _0971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5936__A1 _3983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6783_ _1890_ _1911_ _1912_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4739__A2 net12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8522_ _0085_ _0100_ _0130_ _0115_ _3683_ _3704_ _3717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5734_ _3882_ _0903_ _0904_ _0905_ _0906_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_17_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8453_ _3627_ _3642_ _3657_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5665_ _0377_ _0838_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8320__I _0506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7404_ _2507_ _2515_ _2547_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4616_ _3822_ _3936_ _3937_ _3938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__6361__A1 _1428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8384_ _3536_ _3538_ _3585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5596_ _0768_ _0769_ _0361_ _0770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_7335_ _2471_ _2472_ _2473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4547_ _3860_ _3870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4911__A2 _4225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7266_ _2270_ _2354_ _2398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4478_ _3758_ _3774_ _3791_ _3800_ _3801_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7861__A1 _3018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6217_ _1371_ _1372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6664__A2 _1798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7197_ _2230_ _2323_ _2324_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6148_ _1167_ _1188_ _1306_ _1307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6079_ _1098_ _1109_ _1240_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8642__D _0098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5927__A1 _1089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6015__I _3890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5854__I _0755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5155__A2 _4078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4902__A2 _4216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7852__A1 _0379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5458__A3 _0632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7852__B2 _2872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5863__B1 _1027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4969__A2 _3326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7907__A2 _2579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6591__A1 _1371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8652__CLK clknet_4_11_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5450_ _4080_ _0390_ _0627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5146__A2 _0326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_4_0_Clock_I clknet_3_2_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4401_ _3542_ _2755_ _2764_ A\[3\]\[6\] _3551_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_4
XANTENNA__6894__A2 _2006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5381_ _0553_ _0557_ _0558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_132_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7120_ _2235_ _2240_ _2241_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4332_ _2805_ net7 _2816_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__8096__A1 _3088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7051_ _2044_ _2057_ _2172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7843__A1 _2981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6002_ _1164_ _1020_ _1019_ _1165_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_113_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7953_ _3013_ _3014_ _3123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4843__I _4056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6904_ _3510_ _0013_ _1951_ _2027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7884_ _0293_ _0298_ _3049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_70_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8020__A1 _3184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6835_ _3864_ _1882_ _1961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5909__A1 _0704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6766_ _3767_ _1894_ _1842_ _1895_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_143_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5717_ _0858_ _0859_ _0856_ _0890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8505_ _3702_ _3703_ _0136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6697_ _1822_ _1828_ _1829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_30_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8436_ _3638_ _3639_ _3640_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5648_ _0345_ _0050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8367_ _3564_ _3566_ _3567_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_117_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5579_ A\[2\]\[5\] _4078_ _3271_ _4077_ _0755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4896__A1 _3510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7318_ _2304_ _2453_ _2454_ _2455_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__8087__A1 _3179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8298_ _3455_ _3479_ _3494_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5623__B _0463_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8637__D _0067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7249_ _2295_ _2294_ _2296_ _2291_ _2293_ _2380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_85_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4648__A1 _3965_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7062__A2 _3861_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8675__CLK clknet_4_5_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4820__A1 _3872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6573__A1 _3531_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7117__A3 _2237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4887__A1 _4070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8078__A1 _3160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6089__B1 _1248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7825__A1 _2983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput8 X[3] net8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7053__A2 _2067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8250__A1 _1099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6800__A2 _3775_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4950_ _0058_ _3871_ _4201_ _4264_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_91_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4811__A1 _4112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8002__A1 _3103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4881_ _3144_ _4196_ _4197_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8553__A2 _3687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6620_ _1753_ _1755_ _1756_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5367__A2 _0536_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6551_ _1651_ _1663_ _1692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_119_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5502_ _0546_ _0583_ _0679_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6482_ _1568_ _1578_ _1626_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8221_ _3405_ _3410_ _3411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5433_ _0590_ _0609_ _0610_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6867__A2 _1990_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6331__A4 _3625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8152_ _3334_ _3335_ _3336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5364_ _4056_ _0541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7103_ _2182_ _2220_ _2222_ _2223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4315_ _2578_ _2599_ _2631_ _2642_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_86_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8083_ _3167_ _3237_ _3259_ _3261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5295_ _4089_ _0473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7034_ B\[1\]\[5\] _2155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8698__CLK clknet_4_12_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8241__A1 _3366_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7044__A2 _2164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7936_ _2871_ _2872_ _3104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7867_ _3029_ _2953_ _3030_ _3031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6818_ _1916_ _1917_ _1943_ _1944_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5358__A2 _0398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7798_ _2945_ _2957_ _2958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_52_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6749_ _4200_ _1746_ _1878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_137_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8419_ _3621_ _0107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4748__I _3917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8480__A1 _3678_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4483__I _3805_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5349__A2 _0425_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7034__I B\[1\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7274__A2 _3873_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5080_ _0260_ _0261_ _0262_ _0263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5285__A1 _0374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4393__I _3456_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5588__A2 _0762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5982_ _1039_ _1144_ _1145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7721_ _0334_ _1999_ _2876_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4933_ _4237_ _4246_ _4247_ _4248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8526__A2 _3668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7652_ _2768_ _2779_ _2804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4864_ _3948_ _3824_ _4179_ _4180_ _4181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_32_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6603_ _1739_ _1740_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7583_ _2732_ _2736_ _2738_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4795_ _3326_ _0029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6534_ _1632_ _1634_ _1676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_20_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6465_ _1522_ _1547_ _1609_ _1610_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5416_ _0411_ _0591_ _0592_ _0531_ _0593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_8204_ _3311_ _3318_ _3393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6396_ _1526_ _1542_ _1543_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_115_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8135_ _3316_ _3317_ _3318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4568__I _2745_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5347_ _0454_ _0522_ _0523_ _0524_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8066_ _3241_ _3243_ _3244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5278_ _4089_ _0456_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5276__A1 _0406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7017_ _4135_ _1882_ _2138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7017__A2 _1882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4517__B _3775_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6776__A1 _1838_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5579__A2 _4078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7919_ _3031_ _3035_ _3085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_19_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8650__D _0092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5200__A1 _3048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6700__A1 _3962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8453__A1 _3627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7008__A2 _2128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5019__A1 _0203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6767__A1 _3931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8560__D _0005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5990__A2 _3293_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7192__A1 _2248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput11 X[6] net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4580_ _3843_ _3851_ _3847_ _3902_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_122_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6250_ _1280_ _1401_ _1335_ _1402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__7495__A2 _2592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5201_ _0379_ _0381_ _0382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_42_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4388__I _3402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6181_ _1198_ _1203_ _1337_ _1338_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5132_ _0313_ _0314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_97_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5258__A1 _0023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5063_ _4263_ _0204_ _0246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5025__A4 _0209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5965_ _0993_ _1044_ _1129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_34_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4851__I _4168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7704_ _2814_ _2855_ _2857_ _2858_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_90_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4916_ _4226_ _4229_ _4231_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8684_ _0077_ clknet_4_12_0_Clock C\[3\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5896_ _1059_ _1060_ _1061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5981__A2 _4159_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7635_ _0230_ _0226_ _2788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4847_ _4153_ _4164_ _4165_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7183__A1 _0220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5733__A2 _0873_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7566_ _2650_ _2681_ _2693_ _2720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4778_ _3985_ _4095_ _4097_ _4098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_101_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6778__I _1903_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6517_ _1658_ _1659_ _1660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_88_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7497_ _2645_ _2646_ _2647_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8522__I2 _0130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6448_ _0031_ _0063_ _1513_ _1593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_84_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5497__A1 _0587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4298__I _2449_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6379_ _3981_ _0339_ _1440_ _1438_ _1527_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_88_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8118_ _3208_ _3297_ _3298_ _3299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8645__D _0101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8049_ _3212_ _3213_ _3113_ _3225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6997__A1 _2042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4472__A2 _3787_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6749__A1 _4200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7410__A2 _3929_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6213__A3 _1250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5972__A2 _0030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6921__A1 _1961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8609__CLK clknet_4_11_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8555__D _0000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6988__A1 _2025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5660__A1 _0753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5767__I _0336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5412__A1 _0026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4671__I _3992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5750_ _0774_ _0016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4766__A3 _3964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4701_ _3913_ _4020_ _4021_ _4022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5681_ _0837_ _0852_ _0853_ _0854_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5176__B1 _0355_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7420_ _2561_ _2563_ _2564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4632_ _3931_ _3952_ _3953_ _3954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4563_ _3882_ _0061_ _3884_ _3885_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7351_ _2479_ _2489_ _2490_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6302_ _1452_ _1333_ _1453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7282_ _2400_ _2414_ _2415_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_85_1428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4494_ _3816_ _3817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6233_ _1356_ _1360_ _1385_ _1386_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_116_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6140__A2 _3636_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6164_ _1182_ _1185_ _1320_ _1321_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5115_ _0296_ _0297_ _0298_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_112_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6095_ _3831_ _0569_ _1255_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5046_ _0222_ _0229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5651__A1 _3871_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5651__B2 _4275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6282__B _1432_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6997_ _2042_ _2059_ _2117_ _2118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4581__I _3229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5948_ _1083_ _1112_ _1113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_55_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8667_ _0122_ clknet_4_15_0_Clock C\[2\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5879_ _0988_ _0993_ _1044_ _1045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_55_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7618_ _2742_ _2743_ _2770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_107_1388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6903__A1 _4117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8598_ _0043_ clknet_4_9_0_Clock B\[1\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7549_ _2664_ _2669_ _2702_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_4_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7459__A2 _2604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6131__A2 _1189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4693__A2 _3769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4756__I _3788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5237__A4 _0034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4491__I _3813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7934__A3 _3023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7698__A2 _1865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_3_4_0_Clock_I clknet_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6370__A2 _0063_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6211__I _1249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4381__A1 _3240_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7870__A2 _2562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4684__A2 _3958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8581__CLK clknet_4_4_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7622__A2 _1980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5633__A1 _0804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6920_ _1974_ _1976_ _2043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6851_ _4076_ _0002_ _1976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5802_ _0970_ _0131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5936__A2 C\[2\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6782_ _1893_ _1910_ _1911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_50_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8521_ _3715_ _3716_ _0140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5733_ _0847_ _0873_ _0872_ _0905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8452_ _3627_ _3642_ _3656_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5664_ _0833_ _0834_ _0837_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_50_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7153__A4 _2275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7403_ _2495_ _2506_ _2546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4615_ _3789_ _3937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_8383_ _3581_ _3582_ _3584_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5595_ _3772_ _0354_ _0769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4546_ _3865_ _3868_ _3869_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7334_ _2397_ _2415_ _2472_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7265_ _2332_ _2339_ _2396_ _2397_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4477_ _3794_ _3796_ _3799_ _3800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_137_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6216_ _3972_ _1371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7196_ _2234_ _2241_ _2323_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_58_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4576__I _3897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4675__A2 _3833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6147_ _1171_ _1187_ _1306_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_57_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6078_ _1238_ _1239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5624__A1 _0792_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5029_ _0203_ _0026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7377__A1 _2490_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6352__A2 _1501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7127__I _2055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4363__A1 _3026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7301__A1 _3971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7852__A2 _0381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5458__A4 _0633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4666__A2 _3987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5863__A1 _3777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4486__I _3808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5863__B2 _3926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_11_0_Clock_I clknet_3_5_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6040__A1 _1199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6591__A2 C\[1\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6343__A2 _1492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4400_ _3531_ _3542_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_103_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5380_ _0554_ _0555_ _0556_ _0557_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_126_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4331_ net1 _2805_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7050_ _2044_ _2057_ _2171_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_4_8_0_Clock_I clknet_3_4_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6001_ _1163_ _1164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4396__I _3488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5606__A1 _0776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7952_ _3119_ _3034_ _3120_ _3121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_94_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6903_ _4117_ _0012_ _1948_ _2026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_110_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7883_ _3047_ _0113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6834_ _1884_ _1885_ _1960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6765_ _1840_ _1894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6582__A2 _1720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8504_ _0110_ _3666_ _3703_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5716_ _0835_ _0836_ _0889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6696_ _1824_ _1825_ _1827_ _1828_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_8435_ _3632_ _3637_ _3639_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5647_ _0814_ _0819_ _0820_ _0821_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8366_ _3513_ _3529_ _3565_ _3566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5578_ _0201_ _0052_ _0753_ _0754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_3_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4896__A2 _0029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7317_ _2307_ _2377_ _2454_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4529_ _3843_ _3851_ _3852_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_105_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8297_ _3441_ _3451_ _3493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6098__A1 _1246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7834__A2 _2943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7248_ _2301_ _2378_ _2379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_132_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4648__A2 _3969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7179_ _2302_ _2303_ _2304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8653__D _0070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8506__I _3674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7062__A3 _1755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6270__A1 _0062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4820__A2 _3122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6022__A1 _1184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6573__A2 _1710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7770__A1 _0896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4584__A1 _3904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4887__A2 _4202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8078__A2 _3166_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6089__A1 _0419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6089__B2 _0468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5836__A1 _0310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput9 X[4] net9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8563__D _0008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8250__A2 _1949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4811__A2 _3604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4880_ _0059_ _3870_ _4196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6013__A1 _3993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5775__I _0467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5367__A3 _0543_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6550_ _1687_ _1689_ _1690_ _1691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5501_ _0588_ _0676_ _0677_ _0678_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6481_ _1561_ _1581_ _1625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8220_ _3406_ _3409_ _3410_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5432_ _4130_ _0529_ _0609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8151_ _3244_ _3246_ _3335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5363_ _4010_ _0539_ _0540_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7102_ _2178_ _2221_ _2222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4314_ _2621_ _2631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5294_ _0460_ _0472_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8082_ _3173_ _3258_ _3259_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5827__A1 _4149_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7033_ _2148_ _2149_ _2153_ _2154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__5015__I _0200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5055__A2 _0151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7935_ _3101_ _3036_ _3102_ _3103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7866_ _0401_ _1252_ _1714_ _1736_ _3030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_51_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6817_ _3889_ _0012_ _1918_ _1943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7797_ _2949_ _2954_ _2956_ _2957_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__5358__A3 _0413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6748_ _1831_ _1875_ _1876_ _1855_ _1830_ _1877_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_91_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7504__A1 _2611_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6679_ _1811_ _1812_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8418_ _3618_ _3620_ _3621_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_100_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8648__D _0090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8349_ _3508_ _3532_ _3548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5818__A1 _4028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5818__B2 _4129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8480__A2 _0094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8642__CLK clknet_4_0_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4764__I B\[1\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7991__A1 _0052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6546__A2 _1596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7743__A1 _2839_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8558__D _0003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7274__A3 _1810_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4493__B1 _3745_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5981_ _4215_ _4159_ _1036_ _1144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7982__A1 _3064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7720_ _2873_ _2874_ _2875_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_64_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4796__A1 _0058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4932_ _4241_ _4244_ _4247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7651_ _2768_ _2779_ _2803_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4863_ _3971_ C\[3\]\[8\] _4180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7734__A1 _2799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6602_ _1700_ _1739_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7582_ _2733_ _2735_ _2736_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4794_ _4113_ _0058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6533_ _3434_ _1671_ _1631_ _1674_ _1675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_119_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6464_ _1544_ _1545_ _1543_ _1609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_1448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8203_ _3311_ _3318_ _3392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5415_ _0440_ _0530_ _0592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6395_ _1541_ _1542_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8665__CLK clknet_4_15_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8134_ _0647_ _1851_ _3317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5346_ _0486_ _0521_ _0523_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_115_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8065_ _3060_ _3138_ _3242_ _3243_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8462__A2 _3790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5277_ _0396_ _0405_ _0455_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_101_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6473__A1 _1555_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7016_ _2074_ _2078_ _2137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_130_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4484__B1 _3380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7973__A1 _3052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6776__A2 _1903_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7918_ _3027_ _2995_ _3084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_58_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8517__A3 _3712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7849_ _3009_ _2956_ _3011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_51_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7725__A1 _0488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4533__B _3855_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5200__A2 _2982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4759__I _4079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7135__I _2185_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6700__A2 _1772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4711__A1 _4031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4475__B1 _3797_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4494__I _3816_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5019__A2 _4227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6767__A2 _1725_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7716__A1 _3037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7192__A2 _2286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput12 X[7] net12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8688__CLK clknet_4_5_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4950__A1 _0058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8141__A1 _0899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4669__I _3990_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5200_ _3048_ _2982_ _0380_ _0381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_100_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6180_ _1194_ _1197_ _1337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_48_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5131_ _2599_ net45 _0312_ B\[2\]\[3\] _0313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_123_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7247__A3 _2377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6455__A1 _1598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5258__A2 _0436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5062_ _0238_ _0241_ _0244_ _0245_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_42_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4466__B1 _2826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7955__A1 _3013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5964_ _0985_ _1127_ _1128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7703_ _2807_ _2778_ _2829_ _2857_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4915_ _4226_ _4229_ _4230_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8683_ _0076_ clknet_4_12_0_Clock C\[3\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5895_ _0028_ _0445_ _1060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7634_ _2787_ _0102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4846_ _4156_ _4163_ _4164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_138_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7183__A2 _0015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5194__A1 _3797_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7565_ _2646_ _2684_ _2716_ _2687_ _2719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__8507__I0 _0096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4777_ _3961_ _3824_ _4096_ _4097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_119_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6516_ C\[3\]\[15\] _0947_ _1659_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7496_ _2529_ _2533_ _2593_ _2646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6447_ _1517_ _1520_ _1592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8522__I3 _0115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6378_ _1524_ _1525_ _1526_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8117_ _3219_ _3234_ _3298_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5329_ _0504_ _0505_ _0506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8048_ _3220_ _3223_ _3224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5203__I _0383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8199__A1 _3301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7946__A1 _3113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6749__A2 _1746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8661__D _0130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8371__A1 _0687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6921__A2 _1963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8123__A1 _0509_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7477__A3 _0185_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4448__B1 _2341_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6988__A2 _2094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7937__A1 _0382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8571__D _0016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5412__A2 _0445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4766__A4 _4085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4700_ _3944_ _4019_ _4021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5680_ _0850_ _0851_ _0853_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5176__A1 _0342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4631_ _3771_ _3953_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5176__B2 _0356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7350_ _2483_ _2488_ _2489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4923__A1 _3997_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4562_ _2727_ _3152_ _3884_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_15_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8114__A1 _3281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6301_ _1284_ _1452_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_128_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7281_ _2409_ _2413_ _2414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4493_ _3815_ _3754_ _3745_ _3756_ _3816_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_144_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6232_ _1363_ _1384_ _1385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_100_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6163_ _3794_ _3796_ _1319_ _1179_ _1320_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_112_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6428__A1 _1038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5114_ _0159_ _0174_ _0297_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6094_ _4168_ _0651_ _1254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_111_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5045_ _0227_ _0228_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5023__I _3488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5651__A2 _0050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7928__A1 _3992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4862__I _4092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6996_ _2043_ _2058_ _2117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5179__B _3990_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6600__A1 _0040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5947_ _1086_ _1111_ _1112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_41_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8666_ _0121_ clknet_4_15_0_Clock C\[2\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5878_ _1011_ _1043_ _1044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_55_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8353__A1 _0481_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7617_ _0897_ _1703_ _2769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4829_ _4050_ _4099_ _4147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8597_ _0042_ clknet_4_3_0_Clock B\[1\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6903__A2 _0012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7548_ _2699_ _2700_ _2701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7479_ _2562_ _0006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6682__A4 _1814_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7092__A1 _3240_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4905__A1 _3794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4381__A2 _3326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6658__A1 _1727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4947__I _3845_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8566__D _0011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5330__A1 _3813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6830__A1 _1944_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5778__I _0186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4682__I _3949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6850_ _1975_ _0002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5801_ _0749_ _0969_ _0970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_62_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6781_ _1895_ _1901_ _1909_ _1910_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_95_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8520_ _0114_ _3687_ _3716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5732_ _0847_ _0871_ _0873_ _0904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__8335__A1 _3493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8451_ _3650_ _3654_ _3655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5663_ _0754_ _0758_ _0836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7402_ _2493_ _2516_ _2543_ _2544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4614_ B\[1\]\[3\] _3781_ _2897_ _3784_ _3936_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_8382_ _3544_ _3545_ _3580_ _3582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5594_ _2889_ _0363_ _0768_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7333_ _2400_ _2414_ _2471_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4545_ _3867_ _3122_ _3868_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5018__I _2889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6649__A1 _3972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7264_ _2334_ _2338_ _2396_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_85_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4476_ _3798_ _3799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6215_ _0981_ _0711_ _1370_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7195_ _2321_ _2241_ _2322_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6146_ _1294_ _1304_ _1305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6077_ _1228_ _1237_ _1238_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_57_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6821__A1 _0980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5028_ _0205_ _0212_ _0213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input10_I X[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5388__A1 _2755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6979_ _2100_ _2101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8649_ _0091_ clknet_4_11_0_Clock C\[1\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4363__A2 _3133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5560__A1 _4061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7301__A2 C\[1\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5863__A2 _3789_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7065__A1 _4214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6982__I _2103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8014__B1 _1701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_15_0_Clock_I clknet_3_7_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5379__A1 _4168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6040__A2 _1202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6591__A3 _0468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6879__A1 _1973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5551__A1 _0636_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4330_ _2786_ _2794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_99_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5303__A1 _0479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4677__I _3934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7843__A3 _3003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6000_ _3916_ _3760_ _1163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I K[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7056__A1 _2963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7951_ _3032_ _3033_ _3120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_54_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6902_ _1956_ _2023_ _2024_ _2025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_78_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7882_ _3043_ _3046_ _3047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_36_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6833_ _1887_ _1957_ _1958_ _1959_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6764_ _1891_ _1852_ _1892_ _1893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6560__C _3759_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8503_ _3692_ _3699_ _3700_ _3686_ _3702_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5715_ _0867_ _0887_ _0888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_52_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5790__A1 _0867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6695_ _4215_ _0001_ _1827_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8434_ _3632_ _3637_ _3638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5646_ _0587_ _0672_ _0451_ _0820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_108_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8365_ _3516_ _3528_ _3565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5542__A1 _4218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5577_ _0207_ _0752_ _0753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5971__I _0980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7316_ _2307_ _2377_ _2453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_85_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4528_ _3847_ _3850_ _3851_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8296_ _3438_ _3490_ _3491_ _3481_ _3435_ _3492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_116_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7247_ _2304_ _2307_ _2377_ _2378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_4459_ _2556_ _3782_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_104_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7178_ _2205_ _2214_ _2303_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6129_ _1147_ _1287_ _1288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6307__I _1457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6270__A2 _3905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5211__I _0391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8547__A1 _3693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6022__A2 _4080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7770__A2 _1814_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4584__A2 _3905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8571__CLK clknet_4_6_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4887__A3 _3856_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6089__A2 _0658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7038__A1 _4089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6261__A2 _1331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6217__I _1371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6013__A2 _3790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7761__A2 _1931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5772__A1 _0940_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5500_ _0595_ _0596_ _0594_ _0677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6480_ _1563_ _1580_ _1624_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5431_ _2717_ _0607_ _0608_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_65_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8150_ _3242_ _3333_ _3241_ _3334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5362_ _0353_ _0539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_86_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7101_ _2182_ _2187_ _2221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_82_1207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7277__A1 _0980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4313_ _2610_ _2362_ _2621_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8081_ _3236_ _3258_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5293_ _0463_ _0465_ _0470_ _0471_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_82_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5827__A2 _0989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7032_ _4150_ _2152_ _2153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_141_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7029__A1 _3854_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6252__A2 _1197_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7934_ _3009_ _2955_ _3023_ _3024_ _3102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_42_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7865_ _0720_ _2771_ _1781_ _0383_ _3029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8594__CLK clknet_4_10_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7201__A1 _1768_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6816_ _1940_ _1922_ _1941_ _1942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7796_ _2955_ _2956_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7752__A2 _0012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5358__A4 _0533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5763__A1 _0914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6747_ _1832_ _1854_ _1876_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6678_ _1810_ _1811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5629_ _0792_ _0799_ _0802_ _0803_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8417_ _3581_ _3619_ _3620_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6712__B1 _1842_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8348_ _3512_ _3530_ _3547_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8279_ _0037_ _3302_ _3474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5818__A2 _0982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6779__B1 _1904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7440__A1 _2542_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7991__A2 _1865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4557__A2 _3879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5506__A1 _0606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5809__A2 _0973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7274__A4 _2404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5285__A3 _0462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4493__B2 _3756_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7431__A1 _2510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7431__B2 _2509_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5980_ _1141_ _1142_ _1143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4931_ _4245_ _4246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4796__A2 _0029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7650_ _2798_ _2801_ _2802_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4862_ _4092_ _4179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7734__A2 _2846_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6601_ _1719_ _1730_ _1737_ _1738_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_20_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5745__A1 _0867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7581_ _0920_ _1772_ _2734_ _2735_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4793_ _4112_ _4113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6532_ _3434_ _1671_ _1673_ _1631_ _1674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_101_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6463_ _1594_ _1607_ _1608_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8202_ _3305_ _3306_ _3389_ _3390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5414_ _0590_ _0591_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6394_ _1527_ _1540_ _1541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_115_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8133_ _3312_ _3313_ _3314_ _3316_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5345_ _0486_ _0521_ _0522_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_86_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5026__I _3904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8064_ _3062_ _3137_ _3242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5276_ _0406_ _0373_ _0426_ _0454_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_29_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7015_ _2065_ _2066_ _2136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4865__I _4092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4484__A1 B\[1\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4484__B2 _3756_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6776__A3 _1904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7917_ _3000_ _3082_ _3083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5696__I _0868_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7848_ _3009_ _2956_ _3010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7725__A2 _2771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7779_ _2875_ _2876_ _2936_ _2937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5200__A3 _0380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7489__A1 _2542_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8659__D _0128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7416__I _2502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4711__A2 _3863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4475__A1 B\[1\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4475__B2 _3784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7413__A1 _2498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4778__A2 _4095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7716__A2 _1731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput13 Z[0] net13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8569__D _0014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4950__A2 _3871_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8141__A2 _2614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6152__A1 _4173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5130_ _0305_ _0312_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_97_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5061_ _0239_ _0243_ _0244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4466__A1 A\[2\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4466__B2 _3788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6207__A2 _1265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7955__A2 _3014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5963_ _0973_ _0987_ _1127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4914_ _4228_ _3662_ _4229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_55_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7702_ _2807_ _2778_ _2829_ _2855_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5894_ _0731_ _0734_ _1058_ _1059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8682_ _0075_ clknet_4_11_0_Clock C\[3\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4845_ _4160_ _4162_ _4163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7633_ _2782_ _2785_ _2787_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__7183__A3 _2211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7564_ _2718_ _0093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4776_ _3980_ _4096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8632__CLK clknet_4_11_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8507__I1 _0111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6515_ _1600_ _1657_ _1658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7495_ _2588_ _2592_ _2645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8132__A2 _1894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6446_ _1512_ _1521_ _1591_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6377_ _3999_ _0023_ _1442_ _1525_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
Xclkbuf_4_12_0_Clock clknet_3_6_0_Clock clknet_4_12_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_115_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8116_ _3219_ _3234_ _3297_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5328_ _2755_ _3562_ _0380_ _0505_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_103_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4595__I _3916_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8047_ _3221_ _3222_ _3223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_76_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5259_ _0315_ _0051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4457__A1 _3402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7946__A2 _3114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8371__A2 _2103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8530__I _3724_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5185__A2 _0361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4932__A2 _4244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8123__A2 _1899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7477__A4 _2552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4448__B2 _3770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7937__A2 _0509_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6225__I _0716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8655__CLK clknet_4_12_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4630_ _3761_ _3952_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5176__A2 _0345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4561_ _3883_ _0061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4923__A2 _3818_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8114__A2 _3294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6300_ _1406_ _1450_ _1451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7280_ _2411_ _2412_ _2413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4492_ B\[1\]\[3\] _3815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6231_ _1365_ _1383_ _1384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_48_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6162_ _4182_ _1319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5113_ _0289_ _0294_ _0295_ _0296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6428__A2 _0039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6093_ _0541_ _0037_ _1253_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5044_ _0218_ _0226_ _0227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7928__A2 _0307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8050__A1 _0456_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5939__A1 _1102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6995_ _2035_ _2036_ _2115_ _2116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6600__A2 _1736_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5946_ _1093_ _1110_ _1111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_90_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8665_ _0120_ clknet_4_15_0_Clock C\[2\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5877_ _1013_ _1042_ _1043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_90_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8353__A2 _0007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4828_ _4124_ _4145_ _4146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7616_ _2744_ _2746_ _2768_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8596_ _0041_ clknet_4_3_0_Clock B\[1\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6903__A3 _1948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7547_ _2672_ _2676_ _2700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4759_ _4079_ _4080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8105__A2 _3284_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7478_ _2625_ _2626_ _2627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6429_ _1573_ _1574_ _1575_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_136_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7616__A1 _2744_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7092__A2 _2126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8672__D _0072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8678__CLK clknet_4_7_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7919__A2 _3035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8041__A1 _3210_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6107__A1 _1242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7855__A1 _0514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5330__A2 _0506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5124__I _0305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8280__A1 _0384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8582__D _0027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4841__A1 _4158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8032__A1 _3204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5800_ _0821_ _0968_ _0969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6780_ _1906_ _1908_ _1909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5731_ _0493_ _0903_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5662_ _0833_ _0834_ _0835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_30_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8450_ _3651_ _3652_ _3653_ _3654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7401_ _2490_ _2517_ _2543_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4613_ _3813_ _3934_ _3935_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8381_ _3544_ _3545_ _3580_ _3581_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5593_ _0764_ _0765_ _0766_ _0767_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7332_ _2392_ _2448_ _2468_ _2469_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4544_ _3866_ _3867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7846__A1 _2994_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7263_ _2343_ _2374_ _2393_ _2395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4475_ B\[1\]\[1\] _3781_ _3797_ _3784_ _3798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7514__I _2501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6214_ _1367_ _1257_ _1368_ _1369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7194_ _2234_ _2321_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6145_ _1146_ _1303_ _1304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8546__S _3695_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6076_ _1232_ _1236_ _1237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5027_ _0201_ _0211_ _0212_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6821__A2 _1761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8023__A1 _3109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5388__A2 _3893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6978_ _2099_ _2100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5929_ _0657_ _1094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8648_ _0090_ clknet_4_11_0_Clock C\[1\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8579_ _0024_ clknet_4_6_0_Clock A\[3\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7852__C _3100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5560__A2 _0539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8667__D _0122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7837__A1 _0326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5863__A3 _4182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8262__A1 _3390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7065__A2 _2185_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4823__A1 _4031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8014__A1 _1184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8014__B2 _0577_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5379__A2 _0392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6328__A1 _3636_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6879__A2 _2003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8577__D _0022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5303__A2 _0480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7056__A2 _1863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8253__A1 _0444_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5067__A1 _0025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7950_ _3032_ _3033_ _3119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_23_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6901_ _1959_ _2005_ _2024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_78_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7881_ _3044_ _3045_ _3046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6832_ net39 _1912_ _1958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6567__A1 _2244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6763_ _1837_ _1843_ _1844_ _1892_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_8502_ _0095_ _3676_ _3700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5714_ _0869_ _0885_ _0886_ _0887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6319__A1 _0031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6694_ _1826_ _0001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8433_ _3634_ _3635_ _3637_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5645_ _0817_ _0818_ _0819_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5029__I _0203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8364_ _3553_ _3563_ _3564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5576_ _0751_ _0752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5542__A2 _0718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4527_ _3848_ _3026_ _2706_ _3849_ _3850_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7315_ _2385_ _2451_ _2452_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_89_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8295_ _3452_ _3480_ _3491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_104_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8492__A1 _3689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7246_ _2316_ _2376_ _2377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4458_ _3780_ _3781_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_132_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7177_ _2207_ _2213_ _2302_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4389_ _3413_ _3423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6128_ _1285_ _1286_ _1287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6059_ _1219_ _1220_ _1221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_2_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6751__C _1827_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6022__A3 _4096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5230__A1 _2717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4887__A4 _3857_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5297__A1 _3304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8235__A1 _3351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6013__A3 _4093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5221__A1 _4213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5430_ _0408_ _0607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4688__I _3766_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5361_ _4130_ _0537_ _0538_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7064__I _2086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4312_ net3 _2610_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7100_ _2187_ _2220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8080_ _3254_ _3256_ _3257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7277__A2 _2101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5292_ _4207_ _0467_ _0464_ _0469_ _0470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7031_ _2150_ _2151_ _2152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_102_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7029__A2 _1777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7013__B _2090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6788__A1 _3229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5312__I _3922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7933_ _3009_ _2956_ _3023_ _3024_ _3101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_55_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6852__B _1895_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5460__A1 _0574_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7864_ _2942_ _2943_ _3027_ _3028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6815_ _1877_ _1913_ _1941_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7201__A2 _2100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7795_ C\[0\]\[5\] _4239_ _2955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6746_ _1832_ _1854_ _1875_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6960__A1 _3926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6677_ _1809_ _1810_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8416_ _3539_ _3541_ _3582_ _3585_ _3619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5628_ _0801_ _0796_ _0802_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6712__A1 _4009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8347_ _3506_ _3546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5559_ _0574_ _0537_ _0736_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8278_ _3465_ _3472_ _3473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7229_ _2269_ _2271_ _2284_ _2356_ _2357_ _2358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_59_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8217__A1 _0720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5222__I _0391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6779__A1 _3767_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6779__B2 _0476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8680__D _0073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7991__A3 _3003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6951__A1 _1985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4301__I _2481_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4493__A2 _3754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8590__D _0035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4930_ _4241_ _4244_ _4245_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_3491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7719__B1 _1847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4861_ _4094_ _4097_ _4177_ _4178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6600_ _0040_ _1736_ _1737_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4792_ _2438_ _4112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7580_ _1598_ C\[0\]\[0\] _1630_ _2734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6942__A1 _3969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6531_ _1672_ _1673_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6462_ _1603_ _1606_ _1607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8201_ _0775_ _2562_ _3307_ _3389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5413_ _0398_ _0320_ _0590_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6393_ _1537_ _1539_ _1540_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_47_1103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5344_ _0492_ _0497_ _0520_ _0521_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_8132_ _0631_ _1894_ _3314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5275_ _0452_ _0453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8063_ _3153_ _3239_ _3241_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_47_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7014_ _2068_ _2133_ _2134_ _2135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8561__CLK clknet_4_10_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4484__A2 _3754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7916_ _3005_ _3082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5984__A2 _1146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5198__B B\[0\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7847_ _2954_ _3009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7778_ _2873_ _2874_ _2936_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6933__A1 _2053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6729_ A\[1\]\[4\] _1860_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5217__I _0397_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8675__D _0082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7661__A2 _2813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5672__A1 _0843_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4778__A3 _4097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6924__A1 _3792_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput14 Z[1] net14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4950__A3 _4201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8141__A3 _3128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6152__A2 _0045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8429__A1 _3555_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4702__A3 _4017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8585__D _0030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8584__CLK clknet_4_4_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7101__A1 _2182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7342__I _2359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5060_ _4196_ _0242_ _0243_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6455__A3 _1596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5663__A1 _0754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4466__A2 _3787_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5415__A1 _0440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5962_ _1126_ _0118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5966__A2 _1044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7701_ _2847_ _2853_ _2854_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4913_ _4227_ _3905_ _4228_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8681_ _0074_ clknet_4_7_0_Clock C\[3\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5893_ _0609_ _1057_ _1058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7632_ _2783_ _2784_ _2785_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4844_ _0042_ _4161_ _4162_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7563_ _2691_ _2716_ _2718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4775_ _4086_ _4094_ _4095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8507__I2 _0081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6514_ _1595_ _1602_ _1657_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7494_ _2641_ _2643_ _2644_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6445_ _1508_ _1550_ _1590_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6376_ _1436_ _1523_ _1524_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8115_ _3278_ _3295_ _3296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5327_ _3542_ _2794_ _0331_ B\[0\]\[6\] _0504_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_130_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8046_ _0487_ _2250_ _3222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5258_ _0023_ _0436_ _0437_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5189_ _0367_ _0368_ _0369_ _0370_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_68_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5406__A1 _0548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7159__A1 _1838_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5709__A2 _0880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6906__A1 _1960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5893__A1 _0609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5391__B _3593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4448__A2 _3769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7937__A3 _3104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6950__B _2072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7570__A1 _1673_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4560_ _3877_ _3883_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4491_ _3813_ _3814_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6230_ _1369_ _1378_ _1382_ _1383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_87_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4687__A2 _4007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6161_ _1316_ _1317_ _1318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5112_ _0285_ _0286_ _0295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6092_ _1252_ _0037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7625__A2 _0184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5043_ _0223_ _0225_ _0226_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_112_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7389__A1 _2385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7928__A3 _2237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8050__A2 C\[0\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5939__A2 _1103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6994_ _0202_ _0013_ _2033_ _2115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_80_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5945_ _1098_ _1109_ _1110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_94_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8664_ _0119_ clknet_4_15_0_Clock C\[2\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5876_ _1034_ _1041_ _1042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7615_ _2733_ _2747_ _2767_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4827_ _4127_ _4144_ _4145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_107_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8595_ _0040_ clknet_4_0_0_Clock B\[1\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7546_ _2658_ _2671_ _2699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4758_ _3819_ _4077_ _4078_ A\[2\]\[4\] _4079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_135_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7477_ C\[1\]\[12\] C\[1\]\[13\] _0185_ _2552_ _2626_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4689_ _3830_ _4010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6428_ _1038_ _0039_ _1574_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7864__A2 _2943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6359_ _1410_ _1448_ _1507_ _1508_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7616__A2 _2746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5627__A1 _0800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8029_ _3106_ _3108_ _3202_ _3203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8041__A2 _3214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6052__A1 _1077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4602__A2 _3923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4366__A1 _2727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4905__A3 _3799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7304__A1 _3917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7855__A2 C\[0\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7607__A2 _0010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8280__A2 _2501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8622__CLK clknet_4_1_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6291__A1 _1436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4841__A2 _4152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7791__A1 _0571_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5730_ _0901_ _0902_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_62_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5661_ _0763_ _0771_ _0834_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_88_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4357__A1 _2805_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7400_ _2540_ _2541_ _2542_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4612_ _3933_ _3754_ _3829_ _3756_ _3934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_8380_ _3577_ _3579_ _3580_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_89_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5592_ _0489_ _0199_ _0345_ _0415_ _0766_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7331_ _2395_ _2447_ _2468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_102_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4543_ B\[3\]\[6\] _2930_ _3562_ _2919_ _3866_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_102_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7262_ _2346_ _2372_ _2393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4474_ _3078_ _3797_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_89_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5857__A1 _0043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6213_ _1246_ _1366_ _1250_ _1368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_143_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7193_ _2245_ _2317_ _2318_ _2320_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7059__B1 _1998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6144_ _1298_ _1302_ _1303_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_112_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5609__A1 _0780_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6075_ _1234_ _1235_ _1236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5026_ _3904_ _0211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6821__A3 _1824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7231__B1 _1983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6977_ _2097_ _2098_ _2099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5388__A3 _0380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7782__B2 _1898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4596__A1 _3917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5928_ _1074_ _1092_ _1093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_94_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8647_ _0089_ clknet_4_10_0_Clock C\[1\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5859_ _3822_ _3824_ _4179_ _4180_ _1025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_103_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4348__A1 _2805_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8578_ _0023_ clknet_4_1_0_Clock A\[2\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7529_ _2678_ _2680_ _2681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_5_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7837__A2 _1823_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7301__A4 _2185_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4520__A1 _2449_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8645__CLK clknet_4_9_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8683__D _0076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4823__A2 _3872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8014__A2 _0326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6328__A2 _0711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7828__A2 _2987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5839__A1 _0397_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4511__A1 _3758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8593__D _0038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5067__A2 _4117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4814__A2 _4129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6900_ _1959_ _2005_ _2023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_78_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7880_ _2839_ _2892_ _2901_ _2964_ _2896_ _3045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_63_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6016__A1 _1178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6831_ net39 _1912_ _1957_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6567__A2 _2265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7764__A1 _2909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6762_ _1843_ _1844_ _1837_ _1891_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_1420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8501_ _0080_ _0125_ _3668_ _3699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5713_ _0883_ _0884_ _0886_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6319__A2 _0054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6693_ _1780_ _1826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8432_ C\[0\]\[15\] _1628_ _3635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5644_ _0453_ _0585_ _0812_ _0818_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_15_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8363_ _3555_ _3561_ _3563_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_129_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5575_ _0313_ _0751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7314_ _2387_ _2450_ _2451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8668__CLK clknet_4_15_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4526_ _2963_ _3849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7819__A2 _2915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8294_ _3452_ _3480_ _3490_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7245_ _2320_ _2375_ _2376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4457_ _3402_ _3779_ _3445_ _2513_ _3780_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_63_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4502__A1 _3820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7176_ _2198_ _2290_ _2300_ _2301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_59_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4388_ _3402_ _3413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6127_ _1143_ _1159_ _1286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6058_ _0029_ _0687_ _1220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5009_ C\[3\]\[2\] _0184_ _0195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6558__A2 _3445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4569__A1 _3890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5230__A2 _0315_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8180__A1 _3286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8678__D _0085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4794__I _4113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4727__C _3963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7994__A1 _0049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_3_7_0_Clock clknet_0_Clock clknet_3_7_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_73_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6549__A2 _1628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7746__A1 _2799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6013__A4 _1027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5221__A2 _0401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8546__I0 _0122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8171__A1 _3278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8588__D _0033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5360_ _0362_ _0537_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4311_ _2589_ _2599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_141_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5291_ _0468_ _0469_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6485__A1 C\[2\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7030_ _3894_ _1733_ _2151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6788__A2 _1811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7932_ _3083_ _3087_ _3098_ _3099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_67_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5460__A2 _0493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7863_ _2939_ _2940_ _3027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_64_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6814_ _1877_ _1913_ _1940_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7794_ _2950_ _2951_ _2953_ _2954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_23_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6745_ _1813_ _1817_ _1856_ _1873_ net36 _1874_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_50_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6676_ _1808_ _1809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8162__A1 _3257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4879__I _4195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8415_ _3588_ _3617_ _3618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5627_ _0800_ _0458_ _0466_ _0801_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_118_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6712__A2 _1841_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8346_ _3489_ _3535_ _3545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5558_ _0731_ _0734_ _0735_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_117_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4509_ _3808_ _3832_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_8277_ _3470_ _3471_ _3472_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5489_ _0661_ _0665_ _0666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_132_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6476__A1 _1400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7673__B1 _2824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7228_ _2274_ _2357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_105_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8217__A2 _1987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7159_ _1838_ _2282_ _2283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_76_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6228__A1 _4161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6779__A2 _1907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7728__A1 _2881_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6951__A2 _1894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4962__A1 _4275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5442__A2 _0618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7719__B2 _1850_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4860_ _3978_ _4091_ _4176_ _4177_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_2791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4791_ _3880_ _4040_ _4110_ _4111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6942__A2 _1726_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6530_ _4087_ _1672_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4953__A1 _0028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6461_ _1604_ _1605_ _1606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8200_ _3320_ _3325_ _3387_ _3388_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5412_ _0026_ _0445_ _0589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6392_ _1538_ _0023_ _1539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8131_ _1672_ _3312_ _3313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5343_ _0502_ _0519_ _0520_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_115_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8447__A2 _3462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6458__A1 _1595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8062_ _3155_ _3238_ _3239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_82_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5274_ _0340_ _0449_ _0452_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_130_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7013_ _2072_ _2061_ _2090_ _2134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7958__A1 _0360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5433__A2 _0609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7915_ _3008_ _3079_ _3080_ _3081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7846_ _2994_ _3007_ _3008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_52_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7777_ _2879_ _2885_ _2934_ _2935_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4989_ _0172_ _0173_ _0175_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6933__A2 _2055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6728_ _1859_ _0095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6659_ _1727_ _1729_ _1737_ _1794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8329_ _3520_ _3526_ _3527_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_117_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7110__A2 _2229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5121__A1 _3727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6329__I _1374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5233__I _0413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6773__B _2674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7949__A1 _3023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8691__D _0137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7177__A2 _2213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6999__I _1949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5188__A1 _4169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput15 reset net15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4312__I net3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7101__A2 _2187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5112__A1 _0285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5663__A2 _0758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6612__A1 _3488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5961_ _1120_ _1125_ _1126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_129_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7700_ _2848_ _2852_ _2853_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_59_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4912_ _3888_ _4227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8680_ _0073_ clknet_4_7_0_Clock C\[3\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5892_ _1056_ _1057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5179__A1 _0358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7631_ _2741_ _2752_ _2784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4843_ _4056_ _4161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5718__A3 _0861_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6915__A2 _2037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7562_ _2693_ _2715_ _2716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4926__A1 _4238_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4774_ _4088_ _4091_ _4093_ _3978_ _4094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_105_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6513_ _1604_ _1603_ _1656_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8507__I3 _0126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7493_ _2536_ _2587_ _2643_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6444_ _1589_ _0122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5351__A1 _0492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6375_ _1440_ _1441_ _1523_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8114_ _3281_ _3294_ _3295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5326_ _3315_ _0461_ _0474_ _0503_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8045_ _1252_ _1851_ _3221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5257_ _0435_ _0436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6851__A1 _4076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4457__A3 _3445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5654__A2 _0825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5188_ _4169_ _0360_ _0369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4892__I _4207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5406__A2 _0582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4614__B1 _2897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7159__A2 _2282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7829_ _2979_ _2988_ _2989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_71_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8108__A1 _3186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5228__I _0408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_6_0_Clock clknet_3_3_0_Clock clknet_4_6_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_118_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6768__B A\[0\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8539__I _3731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5893__A2 _1057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7095__A1 _2205_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7937__A4 _2275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4307__I _2383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5138__I _0319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7858__B1 _3020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7781__C _3593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4490_ _3812_ _3813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_144_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5333__A1 _3921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4687__A3 _3805_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6160_ _0044_ _4062_ _1317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5111_ _0285_ _0286_ _0294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_33_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6091_ _0508_ _1252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5042_ _0209_ _0224_ _0225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7302__B _2436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5601__I _0389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6993_ _2039_ _2112_ _2113_ _2114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_92_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5944_ _1100_ _1104_ _1108_ _1109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_55_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8663_ _0118_ clknet_4_14_0_Clock C\[2\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5875_ _1036_ _1040_ _1041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7010__A1 _2064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4826_ _4132_ _4143_ _4144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7614_ _2758_ _2765_ _2766_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8594_ _0039_ clknet_4_10_0_Clock B\[0\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7545_ _2651_ _2696_ _2697_ _2698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4757_ _3787_ _4078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_119_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7476_ _2554_ _2624_ _2625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4688_ _3766_ _4009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_107_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6427_ _1481_ _1572_ _1573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_88_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6358_ _1413_ _1447_ _1507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_66_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7077__A1 _2116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5309_ _0400_ _0487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6289_ _1438_ _1439_ _1440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8028_ _0384_ _1252_ _3104_ _1907_ _3202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_84_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8574__CLK clknet_4_3_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7552__A2 _1630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6760__B1 _1853_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6498__B _1641_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7304__A2 _2350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7855__A3 _0569_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7068__A1 _2174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5660_ _0753_ _0831_ _0832_ _0833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4611_ B\[1\]\[5\] _3933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_90_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5554__A1 _3842_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4357__A2 net6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5591_ _0356_ _0033_ _0765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7330_ _2389_ _2391_ _2467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4542_ _3860_ _3864_ _3865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7261_ _2389_ _2391_ _2392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__7083__I _2126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4473_ _3795_ _3796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5857__A2 _0541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6212_ _1366_ _1250_ _1246_ _1367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7192_ _2248_ _2286_ _2318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7059__A1 _2179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6143_ _1299_ _1301_ _1302_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7059__B2 _3785_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5609__A2 _0782_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6074_ _3905_ _0053_ _0052_ _3899_ _1235_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5025_ _0025_ _0202_ _0205_ _0209_ _0210_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_6_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4293__A1 _2352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6871__B _1995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8597__CLK clknet_4_3_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7231__A1 _1319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7231__B2 _1163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6976_ A\[1\]\[7\] _3709_ _1743_ _2098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_13_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4596__A2 _3814_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5927_ _1089_ _1090_ _1091_ _1092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__6162__I _4182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8646_ _0088_ clknet_4_8_0_Clock C\[1\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5858_ _1022_ _1023_ _1024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_55_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4348__A2 net9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4809_ _4053_ _4125_ _4126_ _4127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_1178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5789_ _0956_ _0957_ _0958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8577_ _0022_ clknet_4_12_0_Clock A\[2\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7528_ _2596_ _2635_ _2679_ _2680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7459_ _2603_ _2604_ _2605_ _2606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4410__I _3636_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5848__A2 _4183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4520__A2 _3842_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4284__A1 B\[3\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8014__A3 _2911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7222__A1 _3817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5536__A1 _4198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7289__A1 _4034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_3_0_Clock clknet_0_Clock clknet_3_3_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__4320__I _2685_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5839__A2 _3863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4511__A2 _3827_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6016__A2 C\[3\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6830_ _1944_ _1955_ _1956_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_36_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6567__A3 _2383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6761_ _4076_ _0001_ _1890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5712_ _0883_ _0884_ _0885_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8500_ _3696_ _3698_ _0135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6692_ _1768_ _1747_ _1825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7516__A2 _0186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5643_ _0815_ _0816_ _0817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8431_ _3601_ _3599_ _3633_ _3634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5527__A1 _4010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8362_ _3559_ _3560_ _3561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5574_ _0750_ _0052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7313_ _2392_ _2448_ _2450_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_116_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4525_ _2889_ _3848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8293_ _3487_ _3489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7244_ _2343_ _2374_ _2375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_85_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4456_ _3727_ _3779_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_85_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7175_ _2201_ _2289_ _2300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_67_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4502__A2 _3822_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4387_ _2233_ _3402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_115_1403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6126_ _1145_ _1158_ _1285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6057_ _1078_ _1217_ _1218_ _1219_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_46_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5008_ _4270_ _0180_ _0194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_2406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6558__A3 _3782_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5766__A1 _0919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4569__A2 _3467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6959_ _3950_ _1971_ _2081_ _2082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_126_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4405__I _2674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8629_ _0103_ clknet_4_8_0_Clock C\[0\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6191__A1 _1232_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8612__CLK clknet_4_2_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8694__D _0140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5297__A3 _0474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6067__I _1089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7994__A2 _2203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8546__I1 _0077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6530__I _4087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4310_ _2319_ net8 _2589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_114_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5290_ _3975_ _0468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8457__I _3660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6485__A2 _1628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7361__I _2282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7434__A1 _0062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7931_ _3090_ _3094_ _3097_ _3098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_83_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5996__A1 _1145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7862_ _3023_ _3024_ _3025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6813_ _1914_ _1921_ _1938_ _1939_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7793_ _0389_ _1894_ _2953_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6744_ _1829_ _1855_ _1873_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4420__A1 _2737_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8635__CLK clknet_4_11_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6675_ _3776_ _1807_ _1808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_104_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5626_ _3845_ _0800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8414_ _3613_ _3616_ _3617_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_30_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5920__A1 _0709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5557_ _0732_ _0733_ _0734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8345_ _3492_ _3534_ _3544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4723__A2 _3953_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4508_ _3830_ _3831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8276_ _0718_ _1987_ _3471_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5488_ _0663_ _0664_ _0665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6476__A2 _1404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7673__A1 _0035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7673__B2 _1534_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7227_ _2280_ _2283_ _2356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4439_ _3761_ _3762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4487__A1 _3806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7158_ _2281_ _2282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6109_ _1227_ _1268_ _1269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_115_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7425__A1 _0061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6228__A2 _0038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7089_ _2175_ _2177_ _2209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_98_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5987__A1 _2685_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7728__A2 _2882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8689__D _0135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4962__A2 _4215_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5911__A1 _0703_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8536__S0 _3678_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7664__A1 _2815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4478__A1 _3758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4478__B2 _3800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7967__A2 _3137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8658__CLK clknet_4_6_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4790_ _4025_ _4039_ _4110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4402__A1 _2330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8599__D _0044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4953__A2 _3889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8144__A2 _3299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6460_ _1526_ _1542_ _1605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5411_ _0214_ _0327_ _0442_ _0447_ _0437_ _0588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_12_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6391_ _3969_ _1538_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8130_ _0514_ C\[0\]\[9\] _3312_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5342_ _0503_ _0511_ _0518_ _0519_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__8447__A3 _0007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8061_ _3167_ _3237_ _3238_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_86_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5273_ _0340_ _0449_ _0450_ _0451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5666__B1 _0775_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7012_ _2072_ _2061_ _2090_ _2133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_29_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7407__A1 _2436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7958__A2 _2077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7914_ _3012_ _3038_ _3080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4641__A1 _3961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7845_ _2997_ _3006_ _3007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_51_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7776_ _2880_ _2884_ _2934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4988_ _0172_ _0173_ _0174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_71_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6727_ _1804_ _1858_ _1859_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6658_ _1727_ _1786_ _1792_ _1793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_125_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5609_ _0780_ _0782_ _0783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6589_ _1371_ C\[1\]\[1\] _1723_ _1726_ _1727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_118_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8328_ _3524_ _3525_ _3526_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_69_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8259_ _3441_ _3451_ _3452_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_106_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4880__A1 _0059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7949__A2 _3109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_2_0_Clock clknet_3_1_0_Clock clknet_4_2_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__4574__B _3821_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4632__A1 _3931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5188__A2 _0360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6385__A1 _1528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6924__A3 _1807_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6137__A1 _0419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8509__S0 _3704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4871__A1 _4167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6612__A2 _1748_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5960_ _1121_ _1124_ _1125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_93_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4623__A1 C\[3\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4911_ _4224_ _4225_ _4226_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5891_ _3625_ _0750_ _1056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8470__I _3668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7630_ _2748_ _2751_ _2783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5179__A2 _0359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4842_ _4157_ _4159_ _4160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6376__A1 _1436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7561_ _2694_ _2698_ _2714_ _2715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_4773_ _4092_ _4093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6512_ _1594_ _1607_ _1654_ _1655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7492_ _2539_ _2586_ _2641_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6443_ _1585_ _1588_ _1589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6374_ _1512_ _1521_ _1522_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_127_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5351__A2 _0497_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5325_ _0500_ _0482_ _0501_ _0502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8113_ _3286_ _3289_ _3292_ _3294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_103_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5256_ _0434_ _0435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8044_ _0403_ _1987_ _3220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6851__A2 _0002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4457__A4 _2513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5187_ _4071_ _0354_ _0368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4614__A1 B\[1\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4614__B2 _3784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8356__A2 _3523_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7828_ _2980_ _2987_ _2988_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_58_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7759_ _0838_ _2120_ _2915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8108__A2 _3189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8513__C1 _3684_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7867__A1 _3029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5342__A2 _0511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4569__B A\[3\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8292__A1 _3371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4853__A1 _4068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8044__A1 _0403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4605__A1 _3423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6803__I _1929_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7858__A1 _3019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7858__B2 _1181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5333__A2 _0509_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5154__I _0335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5110_ _0278_ _0291_ _0292_ _0293_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_112_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6090_ _1249_ _1250_ _1251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8465__I net13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5041_ _0180_ _0189_ _0224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4844__A1 _0042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8035__A1 _3113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6597__A1 _3078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6992_ _2041_ _2093_ _2113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5943_ _1105_ _1106_ _1107_ _1108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_34_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8662_ _0131_ clknet_4_14_0_Clock C\[2\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5874_ _0042_ _1038_ _1039_ _1040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_33_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7010__A2 _2091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7613_ _2762_ _2763_ _2765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4825_ _4139_ _4142_ _4143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_138_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8593_ _0038_ clknet_4_10_0_Clock B\[0\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7544_ _2655_ _2677_ _2697_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4756_ _3788_ _4077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_105_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7475_ C\[1\]\[13\] _0185_ _2624_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4687_ _3952_ _4007_ _3805_ _4008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_134_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer11_I _3572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6426_ _1570_ _1571_ _1572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6357_ _1406_ _1450_ _1506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5308_ _0455_ _0484_ _0485_ _0486_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6288_ _3993_ _1020_ _4176_ _1437_ _4088_ _1439_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5627__A3 _0466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8027_ _3199_ _3129_ _3200_ _3201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6824__A2 _1949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5239_ _3841_ _0419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4835__A1 _4150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4408__I _3615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6623__I _1758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5012__A1 _0192_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6760__A1 _3962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6760__B2 _1836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8697__D _0143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7068__A2 _2188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8017__A1 _2236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6291__A3 _1441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6579__A1 _1688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5251__A1 _3890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5149__I _0330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4610_ _3931_ _3761_ _3921_ _3932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_129_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5590_ _0423_ _0033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5554__A2 _0409_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4541_ _3863_ _3864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7260_ _1768_ _2390_ _2331_ _2329_ _2313_ _2391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_4472_ A\[2\]\[3\] _3787_ _2897_ _3788_ _3795_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_144_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6211_ _1249_ _1366_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7191_ _2248_ _2286_ _2317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6142_ _1296_ _1300_ _1301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7059__A2 _1823_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6073_ _0607_ _0053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6708__I _1839_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5024_ _0207_ _0208_ _0209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8008__A1 _0413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5490__A1 _0655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4293__A2 _2373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7231__A2 _1791_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6975_ net12 _1861_ _2097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5926_ _1037_ _0403_ _1091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6990__A1 _1960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6990__B2 _2028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8645_ _0101_ clknet_4_9_0_Clock C\[1\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5857_ _0043_ _0541_ _1023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4808_ _4054_ _4048_ _4064_ _4126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8576_ _0021_ clknet_4_1_0_Clock A\[2\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5788_ _0914_ _0915_ _0935_ _0957_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_21_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4898__I _3956_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7527_ _2598_ _2634_ _2679_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4739_ _3423_ net12 _4060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7458_ _2103_ _2570_ _2605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6409_ _1405_ _1456_ _1555_ _1556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7389_ _2385_ _2451_ _2530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_66_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8247__A1 _3377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7222__A2 _2350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8691__CLK clknet_4_5_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5536__A2 _0711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7289__A2 _1808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4511__A3 _3833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7213__A2 _2340_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6760_ _3962_ _1772_ _1888_ _1853_ _1836_ _1889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_91_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6972__A1 _2022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5711_ _0850_ _0851_ _0837_ _0884_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_93_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6691_ _4200_ _1823_ _1824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8430_ _3598_ _3602_ _3633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_rebuffer9_I _3604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5642_ _0759_ _0788_ _0816_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5527__A2 _0401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8361_ _3518_ _2665_ _3560_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5573_ _0320_ _0750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6212__B _1246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7312_ _2395_ _2447_ _2448_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8477__A1 _0124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4524_ _2971_ _3846_ _3847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8292_ _3371_ _3433_ _3487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7243_ _2346_ _2372_ _2374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4455_ _3777_ _3778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_104_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7174_ _2299_ _0100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4386_ _3380_ _3391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_113_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4502__A3 _3824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8564__CLK clknet_4_1_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6125_ _1138_ _1191_ _1283_ _1284_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6056_ _1057_ _1079_ _1218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5463__A1 _0637_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5007_ _4270_ _4271_ _4274_ _0193_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_113_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5766__A2 _0932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6958_ _1178_ C\[1\]\[6\] _2081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4569__A3 _2764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5909_ _0704_ _0705_ _1074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6889_ _2012_ _2013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8628_ _0116_ clknet_4_8_0_Clock C\[0\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8559_ _0004_ clknet_4_8_0_Clock A\[0\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4421__I _3735_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8049__B _3113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5206__A1 _3531_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7128__B _2141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4331__I net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8587__CLK clknet_4_1_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7131__A1 _2138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5693__A1 _0864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7434__A2 _2579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8473__I net14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7930_ _3088_ _3095_ _3096_ _3097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_97_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7861_ _3018_ _3021_ _3017_ _3024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6812_ _1915_ _1920_ _1938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7792_ _0383_ net38 _2951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6945__A1 _1984_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6743_ _1866_ _1806_ _1867_ _1872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4420__A2 _3727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6674_ _2897_ _1742_ _1743_ A\[1\]\[3\] _1807_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_52_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8413_ _3546_ _3576_ _3614_ _3616_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5625_ _4198_ _0462_ _0793_ _0799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__7370__A1 _1295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5337__I _0513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8344_ _3543_ _0105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5556_ _3615_ _0529_ _0733_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5920__A2 _0723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4723__A3 _3957_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4507_ _3828_ _3769_ _3829_ _3770_ _3830_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7122__A1 _2225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8275_ _3466_ _3468_ _3469_ _3470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5487_ _3875_ _0658_ _0662_ _0468_ _0664_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_105_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7226_ _2270_ _2348_ _2354_ _2355_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_132_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7673__A2 _1716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4438_ _3760_ _3761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5684__A1 _0835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4487__A2 _3809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7157_ _2150_ _2151_ _3991_ _2281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4369_ B\[3\]\[1\] _2930_ _3207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6108_ _1239_ _1267_ _1268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7425__A2 _2014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7088_ _0059_ _2120_ _2208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5436__A1 _4173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6039_ _1048_ _1200_ _1201_ _1202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5987__A2 _4135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_21 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5739__A2 _0880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6936__A1 _2043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4962__A3 _4220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8536__S1 _3719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7664__A2 _2773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4478__A2 _3774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8293__I _3487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4402__A2 net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5410_ _0453_ _0585_ _0586_ _0587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6390_ _1532_ _1536_ _1537_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8468__I net13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5341_ _0516_ _0517_ _0518_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7104__A1 _2137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8060_ _3173_ _3236_ _3237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7655__A2 _2778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5272_ _0429_ _0448_ _0450_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5666__A1 _0203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5666__B2 _0774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7011_ _2060_ _2092_ _2131_ _2132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6863__B1 _1987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7407__A2 _2499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5418__A1 _0528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8602__CLK clknet_4_9_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7913_ _3012_ _3038_ _3079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4641__A2 _3962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7844_ _3000_ _3005_ _3006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_110_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7775_ _2925_ _2932_ _2933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4987_ _4252_ _4253_ _4233_ _0173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__6394__A2 _1540_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7591__A1 _0436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6726_ _1760_ _1805_ _1857_ _1858_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_109_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6657_ _0179_ _1791_ _1792_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5608_ _0366_ _0370_ _0781_ _0782_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__7894__A2 _2987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6588_ _1725_ _1726_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8327_ _0038_ _3302_ _3525_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5539_ _0648_ _0716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8258_ _3370_ _3450_ _3451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7646__A2 _0011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7209_ _2053_ _2282_ _2337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8189_ _3189_ _3375_ _3376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4880__A2 _3870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6626__I _1761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6082__A1 _1102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output32_I net32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7582__A1 _2733_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6385__A2 C\[3\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6137__A2 _1295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7334__A1 _2397_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8509__S1 _3679_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8625__CLK clknet_4_2_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4871__A2 _4187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8062__A2 _3238_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4484__C _3701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4623__A2 _3929_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4910_ _3865_ _3884_ _4225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_3291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5890_ _0727_ _0743_ _1054_ _1055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4841_ _4158_ _4152_ _4159_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7560_ _2701_ _2713_ _2714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4772_ B\[1\]\[7\] _3780_ _3893_ _3783_ _4092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_140_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6511_ _1605_ _1603_ _1654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7325__A1 _2457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7491_ _2636_ _2639_ _2640_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6442_ _1500_ _1501_ _1586_ _1587_ _1588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_122_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6373_ _1517_ _1520_ _1521_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8112_ _3287_ _3290_ _3291_ _3292_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_138_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5324_ _0499_ _0475_ _0477_ _0501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_88_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8043_ _3209_ _3216_ _3217_ _3219_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5255_ _0430_ _0431_ _0432_ _0433_ _0434_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5186_ _3845_ _0362_ _0367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7827_ _2985_ _2986_ _2987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_12_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7758_ _2810_ _2912_ _2913_ _2864_ _2914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_11_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6709_ _1840_ _1841_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7689_ _2796_ _2831_ _2841_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__8513__B1 _3669_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8513__C2 _0083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8648__CLK clknet_4_11_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4853__A2 _4170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8044__A2 _1987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6055__A1 _1057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4605__A2 _3926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6091__I _0508_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7858__A2 _1770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5869__A1 _4069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8283__A2 _3461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6294__A1 _1429_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5040_ _0219_ _0222_ _0223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4844__A2 _4161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8035__A2 _3114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6046__A1 _0689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6991_ _2041_ _2093_ _2112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7794__A1 _2950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5942_ _0422_ _0720_ _1107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8661_ _0130_ clknet_4_12_0_Clock C\[2\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5873_ _4160_ _4162_ _1039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7612_ _0945_ _1704_ _0010_ _2757_ _2763_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4824_ _4136_ _4140_ _4141_ _4142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_107_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8592_ _0037_ clknet_4_10_0_Clock B\[0\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7543_ _2655_ _2677_ _2696_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4755_ _3818_ _4076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7474_ _1533_ _1983_ _2557_ _2555_ _2622_ _2623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_4686_ _3757_ _4007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6425_ C\[2\]\[14\] _0185_ _1094_ _3898_ _1571_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6356_ _1409_ _1504_ _1505_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5307_ _0471_ _0483_ _0485_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8274__A2 _2055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6287_ _4066_ _0755_ _4179_ _1437_ _1438_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_142_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8026_ _3127_ _3128_ _3200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_76_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5238_ _0416_ _0369_ _0417_ _0418_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8026__A2 _3128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5169_ _0349_ _0350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_56_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7785__A1 _2938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5260__A2 _0051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4424__I _2265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6760__A2 _1772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4771__A1 _4090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4523__A1 _3844_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8265__A2 _3404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6086__I _0456_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8017__A2 _0308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6579__A2 C\[1\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5251__A2 net5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4334__I _2621_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6200__A1 _1242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5003__A2 _0186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4540_ _3862_ _3863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4762__A1 _4076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4471_ _3793_ _3794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5165__I _0330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6210_ _1254_ _1255_ _1364_ _1365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7190_ _2309_ _2315_ _2316_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_48_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8476__I _3675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6141_ _3874_ _0981_ _1300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6072_ _1057_ _1233_ _1234_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4509__I _3808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5023_ _3488_ _0208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6019__A1 _4045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6019__B2 _1181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6974_ _2096_ _0098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5925_ _0541_ _0488_ _1090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8644_ _0100_ clknet_4_8_0_Clock C\[1\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5856_ _1019_ _1021_ _1022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8192__A1 _3375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4807_ _4054_ _4048_ _4064_ _4125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8575_ _0020_ clknet_4_1_0_Clock A\[2\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5787_ _0935_ _0936_ _0942_ _0954_ _0955_ _0956_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_72_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7526_ _2651_ _2655_ _2677_ _2678_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__4753__A1 _4069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4738_ A\[2\]\[7\] _4059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7457_ _2179_ _2390_ _2604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8495__A2 _3674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4669_ _3990_ _3991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6408_ _1453_ _1454_ _1451_ _1555_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7388_ _2457_ _2462_ _2522_ _2528_ _2529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_118_1210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8247__A2 _3382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6339_ _1477_ _1488_ _1489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_7_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4808__A2 _4048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8009_ _0319_ _2045_ _3181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4419__I _2244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6430__A1 _1375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8183__A1 _0750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7930__A1 _3088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4744__A1 _4053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7749__A1 _2847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6421__A1 _1475_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6972__A2 _2025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5710_ _0870_ _0881_ _0882_ _0883_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6690_ _1700_ _1823_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8174__A1 _3299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5641_ _0785_ _0787_ _0815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4999__I _0184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7921__A1 _3084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8360_ _3556_ _3557_ _3558_ _3559_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5572_ _0675_ _0748_ _0749_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_129_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7311_ _2417_ _2446_ _2447_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_89_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4523_ _3844_ _3845_ _3846_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8477__A2 _3669_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8291_ _3486_ _0104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7242_ _2355_ _2371_ _2372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_89_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4454_ _3776_ _3777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5160__A1 _0309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7173_ _2294_ _2297_ _2299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_131_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4385_ _3358_ _3369_ _3380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6124_ _1140_ _1190_ _1283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6055_ _1057_ _1079_ _1217_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6660__A1 _1727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5463__A2 _0638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5006_ _0058_ _3882_ _0192_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5215__A2 _0394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6957_ _2079_ _2000_ _1991_ _2080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_78_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5908_ _0735_ _0741_ _1072_ _1073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8165__A1 _3262_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6888_ _2011_ _2012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5839_ _0397_ _3863_ _1005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8627_ _0115_ clknet_4_8_0_Clock C\[0\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7912__A1 _3064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4726__A1 _3993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8558_ _0003_ clknet_4_8_0_Clock A\[0\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7509_ _2100_ _2616_ _2659_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8489_ _3685_ _3688_ _0133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7140__A2 _2261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5151__A1 _3892_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5151__B2 B\[0\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5533__I _0656_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5206__A2 _2786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6167__B1 _1322_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7903__A1 _2981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5390__A1 _3978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8459__A2 _3799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5142__A1 _0309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7434__A3 _2402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7860_ _3022_ _3023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_91_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6811_ _1815_ _1935_ _1936_ _1937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_93_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7791_ _0571_ _1714_ _2950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6945__A2 _2067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6742_ _1805_ _1868_ _1869_ _1858_ _1870_ _1800_ _1871_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai33_1
XFILLER_108_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8147__A1 _3257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4420__A3 _2373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6673_ _1765_ _0010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4522__I _2695_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5624_ _0792_ _0797_ _0798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4708__A1 _3846_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8412_ _3549_ _3575_ _3614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7370__A2 _1949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8343_ _3539_ _3541_ _3543_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5555_ _3304_ _0319_ _0732_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4506_ _3185_ net10 _3829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8274_ _0631_ _2055_ _3469_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5486_ _3133_ _0657_ _0662_ _0663_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__7122__A2 _2242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7225_ _2349_ _2351_ _2353_ _2354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_132_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4437_ _3759_ _3760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_104_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8681__CLK clknet_4_7_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7156_ _2277_ _2279_ _2280_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4368_ _3185_ net6 _3196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_116_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6107_ _1242_ _1266_ _1267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7087_ _2174_ _2188_ _2206_ _2207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4299_ net1 _2470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_1470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5436__A2 _4026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6038_ _0972_ _1046_ _1201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7189__A2 _2314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5739__A3 _0870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6936__A2 _2058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7989_ _3087_ _3098_ _3159_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_1537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7664__A3 _1771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6872__A1 _3802_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6624__A1 _3904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4607__I _3928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8129__A1 _3309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8554__CLK clknet_4_14_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4342__I _2908_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5363__A1 _4010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6560__B1 _1699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5340_ _0512_ _0466_ _0515_ _3976_ _0517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8301__A1 _3378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6269__I _3874_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5271_ _0429_ _0448_ _0449_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_49_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5173__I _0353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7010_ _2064_ _2091_ _2131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5666__A2 _0838_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6863__A1 _1985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6863__B2 _4012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7912_ _3064_ _3076_ _3077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_48_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8368__A1 _3497_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4641__A3 _3796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7843_ _2981_ _3001_ _3003_ _3005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_93_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4986_ _0161_ _0170_ _0171_ _0172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7774_ _2926_ _2931_ _2932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_75_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7591__A2 _1826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6725_ _1806_ _1818_ _1856_ _1857_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_6656_ net34 _1791_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8540__A1 _0091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7343__A2 _2428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5607_ _0309_ _0316_ _0321_ _0781_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__5354__A1 _0310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6587_ _1724_ _1725_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5538_ _0713_ _0714_ _0715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8326_ _3521_ _3522_ _3523_ _3524_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8257_ _3444_ _3449_ _3450_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5469_ _0568_ _0646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7208_ _4133_ _1809_ _2336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8188_ _3992_ _0576_ _3002_ _3375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_114_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7139_ _4035_ _1746_ _2261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6606__A1 _3358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6082__A2 _1103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4427__I _3749_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8359__A1 _3462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4632__A3 _3953_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8577__CLK clknet_4_12_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6909__A2 _2031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6642__I _1710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7582__A2 _2735_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6385__A3 A\[2\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7473__I _2498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5896__A2 _1060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7098__A1 _2135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4337__I _2856_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7270__A1 _3864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4623__A3 _3939_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7022__A1 _2137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4840_ _4066_ _4158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5584__A1 _0754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4771_ _4090_ C\[3\]\[7\] _4091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6510_ _1512_ _1521_ _1611_ _1652_ _1653_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_7490_ _2637_ _2638_ _2639_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7325__A2 _2462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6441_ _1458_ _1460_ _1499_ _1587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6372_ _1300_ _1518_ _1422_ _1519_ _1520_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_31_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8111_ _0409_ _1864_ _3291_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5323_ _0475_ _0477_ _0499_ _0500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8042_ _3215_ _3210_ _3214_ _3217_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5254_ B\[0\]\[0\] _0433_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5185_ _0357_ _0361_ _0365_ _0366_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7013__A1 _2072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7826_ _2759_ _2014_ _2986_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4969_ _4227_ _3326_ _0155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7757_ _0335_ _0752_ _2911_ _1702_ _0761_ _2913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_6708_ _1839_ _1840_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8513__A1 _0113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7316__A2 _2377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7688_ _2796_ _2831_ _2840_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8513__B2 _0128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5327__A1 _3542_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6639_ _1769_ _1773_ _1774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_137_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4710__I _2878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8309_ _3503_ _3505_ _3506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_133_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6637__I _1771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6055__A2 _1079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5566__A1 _0730_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4369__A2 _2930_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8504__A1 _0110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5318__A1 _3773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5869__A2 _0020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6547__I _1598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8035__A3 _3116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7243__A1 _2346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6990_ _1960_ _1969_ _2037_ _2038_ _2028_ _2111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_66_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7794__A2 _2951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5941_ _3805_ _0646_ _1106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8660_ _0129_ clknet_4_14_0_Clock C\[2\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5872_ _1037_ _1038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4823_ _4031_ _3872_ _4141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7611_ _2761_ _0008_ _1759_ _2757_ _2762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_21_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8591_ _0036_ clknet_4_9_0_Clock B\[0\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7542_ _2673_ _2675_ _2694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4754_ _4046_ _4068_ _4074_ _4044_ _4075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7473_ _2498_ _2622_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4685_ _4000_ _4005_ _4006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5626__I _3845_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4530__I _2481_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6424_ _1528_ C\[2\]\[14\] B\[2\]\[7\] _3898_ _1570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_128_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6355_ _1449_ _1504_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7841__I _1807_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5306_ _0471_ _0483_ _0484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_88_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6286_ _0456_ C\[3\]\[12\] _1437_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8025_ _3127_ _3128_ _3199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5237_ _4073_ _4262_ _0414_ _0034_ _0417_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_9_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4835__A3 _4152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5168_ _2610_ _2362_ _0349_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5099_ _0273_ _0282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5796__A1 _0866_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4705__I _3304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7809_ _2967_ _0959_ _2968_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8615__CLK clknet_4_1_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4771__A2 C\[3\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4440__I B\[1\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4523__A2 _3845_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6367__I _1419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4287__A1 _2330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8017__A3 _3002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5236__B1 _0034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7776__A2 _2884_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6579__A3 _1630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4615__I _3789_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4762__A2 _0020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4350__I _2993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4470_ _3792_ _3793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6140_ _3883_ _3636_ _1299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6071_ _3898_ _0607_ _1233_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5181__I _0344_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5475__B1 _0651_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5022_ _0206_ _0207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6019__A2 _4067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6973_ _2016_ _2019_ _2095_ _2096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__4525__I _2889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5924_ _1087_ _0721_ _1088_ _1089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8638__CLK clknet_4_9_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6990__A3 _2037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8643_ _0099_ clknet_4_8_0_Clock C\[1\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5855_ _4001_ _3948_ _1020_ _1021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__8192__A2 _3378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4806_ _3869_ _4037_ _4123_ _4124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8574_ _0019_ clknet_4_3_0_Clock A\[2\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5786_ _0919_ _0932_ _0942_ _0955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_7525_ _2672_ _2676_ _2677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_120_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4737_ _3955_ _4007_ _3831_ _4058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__4753__A2 _4070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5356__I _0353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4668_ _2663_ _3990_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7456_ _2485_ _2484_ _2603_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6407_ _1552_ _1553_ _1554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5702__A1 _0848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7387_ _2452_ _2455_ _2528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4599_ _3920_ _3921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_116_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6338_ _1484_ _1487_ _1488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_1_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6269_ _3874_ _0062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8008_ _0413_ _2012_ _3180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7207__A1 _3863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6430__A2 _1482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8183__A2 _2101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5941__A1 _3805_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5457__B1 _0633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4432__A1 _3727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6972__A3 _2094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5640_ _0812_ _0813_ _0814_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5571_ _0678_ _0681_ _0747_ _0748_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_79_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4522_ _2695_ _3845_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7310_ _2419_ _2445_ _2446_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_102_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8290_ _3424_ _3485_ _3486_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8487__I _3686_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7241_ _2358_ _2370_ _2371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4453_ _3775_ _3776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7172_ _2295_ _2296_ _2297_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4384_ net5 _3369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_113_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6123_ _1132_ _1133_ _1137_ _1282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7437__A1 _2573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6054_ _1214_ _1215_ _1216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5005_ _0188_ _0190_ _0191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6660__A2 _1729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6735__I _1865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6956_ _4003_ _1770_ _1990_ _4088_ _2079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5907_ _1070_ _1071_ _0740_ _1072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_22_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6887_ _2010_ _3776_ _1861_ _1698_ _3967_ _2011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_70_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8602__D _0047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8626_ _0114_ clknet_4_2_0_Clock C\[0\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5838_ _3868_ _1002_ _1003_ _4140_ _1004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_33_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8557_ _0002_ clknet_4_2_0_Clock A\[0\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5923__A1 _4218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5769_ _0927_ _0938_ _0939_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_124_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7508_ _2656_ _2657_ _2658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8488_ _0068_ _3687_ _3669_ _0070_ _3688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7439_ _2544_ _2584_ _2585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5814__I _3026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5151__A2 _3391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6100__A1 _1105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6645__I _1779_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4662__A1 _3983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5206__A3 _0330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6380__I _1372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6167__A1 _3961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6167__B2 _4088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7903__A2 _3003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4717__A2 _4037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5914__A1 _3897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5390__A2 _0566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7667__A1 _0924_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5724__I _0343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7419__A1 _1538_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8092__A1 _3262_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6810_ net35 _1923_ _1936_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7790_ C\[0\]\[4\] _3929_ _2938_ _2948_ _2949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_51_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6741_ _1722_ _1751_ _1870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4956__A2 _3922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8147__A2 _3261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6158__A1 _0045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6672_ _1767_ _1798_ _1806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8411_ _3589_ _3610_ _3612_ _3613_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_5623_ _0794_ _0796_ _0463_ _0797_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4708__A2 _4028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8342_ _3424_ _3485_ _3540_ _3541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5554_ _3842_ _0409_ _0731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7658__A1 _0050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4505_ A\[2\]\[5\] _3828_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5485_ _3972_ C\[2\]\[8\] _0662_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8273_ _1672_ _3466_ _3468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4436_ _3691_ _3759_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7224_ _3969_ _0003_ _2353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6330__A1 _1479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4367_ _2330_ _3185_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7155_ _1018_ _2275_ _2278_ _2279_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_98_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6106_ _1259_ _1265_ _1266_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7086_ _2173_ _2189_ _2206_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4298_ _2449_ _2460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7830__A1 _2879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5436__A3 _0364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6037_ _0972_ _1046_ _1200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6397__A1 _1433_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7988_ _3156_ _3157_ _3158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6939_ _1989_ _2001_ _2062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_78 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6149__A1 _0021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8609_ _0054_ clknet_4_11_0_Clock B\[2\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5372__A2 _0495_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7649__A1 _2799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8310__A2 _3505_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6321__A1 _0327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7664__A4 _1972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6872__A2 _1710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4883__A1 _2460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6624__A2 _1740_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6388__A1 _1479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5060__A1 _4196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6560__A1 _3380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5363__A2 _0539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6560__B2 A\[1\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5454__I _0630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8301__A2 _3496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5270_ _0437_ _0447_ _0448_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_99_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6863__A2 _1783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7812__A1 _2904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7911_ _3066_ _3075_ _3076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_55_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7842_ _3793_ _0751_ _3002_ _3003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__6379__A1 _3981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7040__A2 _2159_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7773_ _2927_ _2929_ _2931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4929__A2 _3923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4985_ _0168_ _0169_ _0171_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6724_ _1821_ _1830_ _1855_ _1856_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_108_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6655_ _1788_ _1789_ _3759_ _1790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8540__A2 _3676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5606_ _0776_ _0779_ _0780_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5354__A2 _0408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6586_ _3759_ _1708_ _1712_ _1724_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_118_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8325_ _0631_ _2087_ _3523_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5537_ _4198_ _0711_ _0712_ _0469_ _0714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5364__I _4056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8256_ _3447_ _3448_ _3449_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5468_ _0642_ _0643_ _0644_ _0645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7207_ _3863_ _2045_ _2335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5657__A3 _0765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4419_ _2244_ _3727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_8_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8187_ _1099_ _1765_ _1810_ _0444_ _3374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5399_ _3894_ _0304_ _0306_ B\[2\]\[7\] _0576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_119_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7138_ _2258_ _2259_ _2260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_86_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6409__B _1555_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7803__A1 _2904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7069_ _2173_ net40 _2190_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_86_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4617__A1 _3932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8359__A2 _0006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7031__A2 _2151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5042__A1 _0209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5539__I _0648_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6385__A4 _0047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5593__A2 _0765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7098__A2 _2170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8295__A1 _3452_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4608__A1 C\[3\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7270__A2 _1928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5820__A3 _0984_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4353__I _2737_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5584__A2 _0758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6781__A1 _1895_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4770_ _4089_ _4090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8671__CLK clknet_4_4_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8700__D _0146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6440_ _1458_ _1460_ _1499_ _1586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6533__A1 _3434_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6371_ _1420_ _1513_ _1519_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_115_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8110_ _0443_ _1809_ _3290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5322_ _0419_ _0498_ _0464_ _0499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8041_ _3210_ _3214_ _3215_ _3216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5253_ _3413_ _3467_ _0380_ _0432_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_87_106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4847__A1 _4153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8038__A1 _0718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5184_ _0356_ _3848_ _0364_ _0355_ _0365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_69_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7261__A2 _2391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8210__A1 _1181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7825_ _2983_ _2984_ _2985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_52_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5024__A1 _0207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7756_ _4158_ _0761_ _2911_ _2912_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_51_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4968_ _0152_ _0153_ _0154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6707_ _1790_ _1839_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_138_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7687_ _2792_ _2833_ _2838_ _2839_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_4899_ _3757_ _4214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8513__A2 _3708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5327__A2 _2794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6638_ _3786_ _1772_ _1773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6569_ _3358_ _3369_ _1707_ _1708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8308_ _3444_ _3449_ _3504_ _3505_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6288__B1 _1437_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8239_ _3359_ _3416_ _3429_ _3430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6827__A2 _1952_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8029__A1 _3106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4438__I _3760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7252__A2 _2314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8694__CLK clknet_4_7_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8201__A1 _0775_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4774__B1 _4093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8504__A2 _3666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5318__A2 _0401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5869__A3 _4068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6563__I _1702_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5940_ _4072_ _0649_ _1105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5871_ _4062_ _1037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5006__A1 _0058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7610_ _2760_ _2761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4822_ _2685_ _3862_ _4140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8590_ _0035_ clknet_4_2_0_Clock B\[0\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6754__A1 _4202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7541_ _2678_ _2692_ _2693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4753_ _4069_ _4070_ _4073_ _4074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7472_ _2612_ _2619_ _2620_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4684_ _3918_ _3958_ _4004_ _3938_ _4005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_135_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6423_ _1485_ _1486_ _1569_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_105_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8259__A1 _3441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6354_ _1503_ _0121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5305_ _0465_ _0478_ _0482_ _0483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__8567__CLK clknet_4_0_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6285_ _1324_ _1326_ _1435_ _1436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_3_0_Clock_I clknet_3_1_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8024_ _3168_ _3195_ _3197_ _3169_ _3170_ _3198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_130_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5236_ _4262_ _0414_ _0034_ _4073_ _0416_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5167_ _0347_ _0348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_5_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5098_ _0247_ _0279_ _0280_ _0281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7785__A3 _2943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8605__D _0050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5796__A2 _0964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7808_ _0934_ _0958_ _2967_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7739_ _2894_ _0081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8498__A1 _3679_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4287__A2 net7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7479__I _2562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5236__B2 _4073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7933__B1 _3023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6332__B _1481_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5727__I _0823_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4631__I _3771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7942__I C\[0\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6070_ _1229_ _1230_ _1231_ _1092_ _1074_ _1232_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_112_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5475__A1 _3772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input9_I X[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5021_ _4033_ _0206_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5475__B2 _3956_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6019__A3 _4093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6972_ _2022_ _2025_ _2094_ _2095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_47_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6975__A1 net12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5923_ _4218_ _4273_ _0647_ _0649_ _1088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8642_ _0098_ clknet_4_0_0_Clock C\[1\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5854_ _0755_ _1020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4805_ _4030_ _4038_ _4123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8573_ _0018_ clknet_4_3_0_Clock A\[2\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5785_ _0941_ _0953_ _0954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4541__I _3863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7524_ _2673_ _2675_ _2676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_72_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4736_ _3955_ _4009_ _4056_ _4057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_119_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4753__A3 _4073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7455_ _2600_ _2601_ _2602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4667_ _3758_ _3827_ _3989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_107_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6406_ _1505_ _1506_ _1551_ _1553_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_116_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7386_ _2527_ _0089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4598_ _3919_ _3744_ _3196_ _3750_ _3920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_66_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6337_ _1485_ _1486_ _1487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_103_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6268_ _3326_ _1419_ _1420_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8007_ _3121_ _3131_ _3178_ _3179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_9_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5219_ _0379_ _0381_ _3946_ _0400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_76_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6199_ _1221_ _1349_ _1353_ _1354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_28_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8404__A1 _3555_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7207__A2 _2045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5218__A1 _0398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6966__A1 _2080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6931__I _1998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4744__A3 _4064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7694__A2 _0011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7446__A2 _2592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5457__A1 _3965_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5457__B2 _4213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5209__A1 _3701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4626__I _3947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7002__I _2013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8542__B _3708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4432__A2 _2373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4361__I _3111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5570_ _0693_ _0746_ _0747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_129_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4521_ _3015_ _3844_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7240_ _2361_ _2369_ _2370_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4452_ _2856_ _3775_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_144_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7171_ _2016_ _2104_ _2110_ _2194_ _2105_ _2296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_4383_ _2319_ _3358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6122_ _1128_ _1279_ _1280_ _1281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6053_ _1073_ _1082_ _1215_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5999__A2 _1041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5004_ _0180_ _0189_ _0190_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8605__CLK clknet_4_0_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4536__I _3858_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6955_ _3832_ _2077_ _2078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5620__A1 _0342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7847__I _2954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5906_ _0736_ _0737_ _1071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6886_ A\[1\]\[6\] _2010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8625_ _0113_ clknet_4_2_0_Clock C\[0\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5837_ _4136_ _4141_ _1003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7373__A1 _2510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8556_ _0001_ clknet_4_2_0_Clock A\[0\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5768_ _0016_ _0925_ _0938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4726__A3 _3950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5923__A2 _4273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7507_ _2620_ _2630_ _2657_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4719_ _4025_ _4039_ _4040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_5_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8487_ _3686_ _3687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7125__A1 _2147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5699_ _0871_ _0872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7438_ _2569_ _2583_ _2584_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_107_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7369_ _2440_ _2441_ _2510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_89_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5151__A3 _0331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5439__A1 _4056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6100__A2 _1106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4662__A2 C\[3\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4446__I _3735_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6939__A1 _1989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5611__A1 _0773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7364__A1 _2502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6167__A2 _4079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5914__A2 _0051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7667__A2 _1975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8628__CLK clknet_4_8_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7419__A2 _2562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6836__I _1902_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4356__I _2786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5602__A1 _0774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6571__I _1709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6740_ _1760_ _1857_ _1869_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4956__A3 _3767_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6671_ _1801_ _1799_ _1805_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6158__A2 _4161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8410_ _3567_ _3574_ _3611_ _3612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5622_ _0795_ _0458_ _0466_ _2717_ _0796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_125_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8341_ _3427_ _3484_ _3540_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7107__A1 _3015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5553_ _0629_ _0728_ _0729_ _0730_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4504_ _3709_ _3766_ _3804_ _3827_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_121_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8272_ _0457_ C\[0\]\[11\] _3466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7658__A2 _1762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5484_ _0575_ _0659_ _0660_ _0661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5669__A1 _3973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7223_ _1962_ _0003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4435_ _3709_ _3751_ _3757_ _3758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__6330__A2 C\[2\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7154_ _0513_ C\[1\]\[8\] _2652_ _2278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4366_ _2727_ _3152_ _3163_ _3174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6618__B1 _1743_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6105_ _1262_ _1264_ _1265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_141_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5650__I _0822_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7085_ _2202_ _2204_ _2205_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4297_ _2438_ _2449_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6094__A1 _4168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6036_ _4261_ _0178_ _0300_ _1047_ _1199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5436__A4 _0355_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5841__A1 _1002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6397__A2 _1443_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7987_ _2760_ _2103_ _3073_ _3157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7594__A1 _2744_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_35 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8613__D _0058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6938_ _1989_ _2001_ _2061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6869_ _1991_ _1993_ _1994_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7346__A1 _3874_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6149__A2 _3999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8608_ _0053_ clknet_4_11_0_Clock B\[2\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5357__B1 _0533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7897__A2 _3039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8539_ _3731_ _0145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4332__A1 _2805_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4885__B _3794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4883__A2 _4198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6656__I net34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6085__A1 _0374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7821__A2 _2932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5832__A1 _4153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7585__A1 _0209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6388__A2 C\[3\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6391__I _3969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6560__A2 _1698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4571__A1 _3358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4323__A1 _2460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6566__I _3809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6076__A1 _1232_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7273__B1 _2404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5823__A1 _4165_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7910_ _3073_ _3074_ _3075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_95_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7841_ _1807_ _3002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_24_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7576__A1 _2721_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6379__A2 _0339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7772_ _2912_ _2928_ _2929_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4984_ _0168_ _0169_ _0170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_52_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6723_ _1831_ _1832_ _1854_ _1855_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__7328__A1 _2387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6654_ _2341_ _1710_ _1789_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6000__A1 _3916_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5605_ _0777_ _0778_ _0394_ _0779_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_30_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6585_ B\[1\]\[1\] _1723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8324_ _1672_ _3521_ _3522_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4562__A1 _2727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5536_ _4198_ _0711_ _0712_ _0713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_121_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8255_ _0607_ _2123_ _3448_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5467_ _0560_ _0580_ _0644_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7860__I _3022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7206_ _2235_ _2240_ _2333_ _2334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4418_ A\[2\]\[3\] _3718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8186_ _3371_ _3372_ _3373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5398_ _0574_ _0472_ _0575_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7137_ _3968_ _1841_ _2259_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8608__D _0053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4349_ _2982_ _2908_ _2298_ B\[3\]\[4\] _2993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7068_ _2174_ _2188_ _2189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6606__A3 _2373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4617__A2 _3935_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6019_ _4045_ _4067_ _4093_ _1179_ _1181_ _1182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_27_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4724__I _3947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7100__I _2187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6058__A1 _0029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4608__A2 _3826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7558__A1 _2659_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4634__I _3920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8550__B _3675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5465__I _0573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7730__A1 _2879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6533__A2 _1671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6370_ _3646_ _0063_ _1518_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5321_ _0461_ _0498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8040_ _3018_ _3215_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_3_3_0_Clock_I clknet_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5252_ _3892_ _0331_ _0431_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8038__A2 _1736_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5183_ _0363_ _0364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_64_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7824_ _0838_ _1952_ _2984_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5024__A2 _0208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7755_ _1744_ _2911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4967_ _4199_ _4204_ _0153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6706_ _3766_ _1838_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7686_ _2783_ _2782_ _2832_ _2838_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4898_ _3956_ _4213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6637_ _1771_ _1772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7721__A1 _0334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5327__A3 _0331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4535__A1 _3760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6568_ _1706_ _1707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_4_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5519_ _0645_ _0667_ _0696_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8307_ _3370_ _3450_ _3504_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6499_ _1624_ _1625_ _1641_ _1643_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__6288__A1 _3993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8238_ _3362_ _3415_ _3429_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6288__B2 _4088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmultiply_komal_33 done vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_105_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8169_ _3352_ _3353_ _3354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7788__A1 _0387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6460__A1 _1526_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5263__A2 _0440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4454__I _3776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8201__A2 _2562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4774__A1 _4088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4774__B2 _3978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7005__I _2102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6451__A1 _4152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4462__B1 _2826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5870_ _4171_ _4174_ _1035_ _1036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5006__A2 _3882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_10_0_Clock_I clknet_3_5_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4821_ _4134_ _4136_ _4138_ _4032_ _4139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XTAP_2390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6754__A2 _1882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7540_ _2680_ _2692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4752_ _4072_ _4073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4765__B2 _3765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7471_ _2616_ _2618_ _2619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5195__I _0375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4683_ _4001_ _3778_ _4002_ _4003_ _3979_ _4004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__4517__A1 _3838_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6422_ _1566_ _1567_ _1568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5190__A1 _0366_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6353_ _1461_ _1499_ _1502_ _1503_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__8259__A2 _3451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5304_ _3997_ _0481_ _0482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6284_ _1184_ _4080_ _4176_ _1322_ _1435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_130_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8023_ _3109_ _3117_ _3197_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4539__I _3861_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5235_ _0415_ _0034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5166_ _2492_ _3782_ _0346_ B\[0\]\[2\] _0347_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_57_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_7_0_Clock_I clknet_3_3_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5097_ _0263_ _0274_ _0280_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8195__A1 _3377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7807_ _2966_ _0082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5999_ _1034_ _1041_ _1161_ _1162_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8621__D _0102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7738_ _0259_ _0275_ _0256_ _2894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_138_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8498__A2 _3678_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7669_ _2820_ _2821_ _2822_ _2823_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_14_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4449__I _3771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8661__CLK clknet_4_12_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5236__A2 _0414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8186__A1 _3371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4912__I _3888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4747__A1 _4066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5172__A1 _0348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4359__I _2856_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5020_ _0204_ _0205_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5475__A2 _0569_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4683__B1 _4003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6424__A1 _1528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6971_ _2039_ _2041_ _2093_ _2094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_80_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5922_ _4218_ _0647_ _0649_ _3773_ _1087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_59_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8641_ _0097_ clknet_4_0_0_Clock C\[1\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5853_ _3761_ _4168_ _1018_ _1019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_61_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7924__A1 _0363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4804_ _4041_ _4101_ _4121_ _4122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5784_ _0944_ _0952_ _0953_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8572_ _0017_ clknet_4_3_0_Clock A\[2\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7523_ _2570_ _2604_ _2675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4735_ _4014_ _4056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7454_ _2574_ _2565_ _2601_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4666_ _3945_ _3987_ _3988_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_31_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6405_ _1505_ _1506_ _1551_ _1552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7385_ _2522_ _2526_ _2527_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4597_ A\[2\]\[1\] _3919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8684__CLK clknet_4_12_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4910__A1 _3865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6336_ _1038_ _0038_ _1486_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6267_ _1295_ _1419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8006_ _3126_ _3130_ _3178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_88_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5218_ _0398_ _0377_ _0399_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6198_ _1352_ _1353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_44_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6484__I _0947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8616__D _0061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5149_ _0330_ _0331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6415__A1 _0327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5218__A2 _0377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6966__A2 _2085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8168__A1 _3270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4729__A1 _4048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4901__A1 _4070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6654__A1 _2341_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5457__A2 _0632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7851__B1 _1732_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5209__A2 _0389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8557__CLK clknet_4_2_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4642__I _3813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7382__A2 _2455_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5393__A1 _3921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4520_ _2449_ _3842_ _3843_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4451_ _3762_ _3767_ _3773_ _3774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_7_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7170_ _2110_ _2194_ _2295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4382_ _3174_ _3337_ _3347_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6121_ _1131_ _1192_ _1280_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6052_ _1077_ _1081_ _1214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5003_ C\[3\]\[0\] _0186_ _0189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4817__I _4034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8398__A1 _1597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7070__A1 _2135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6954_ _2075_ _2076_ _2077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5620__A2 _0498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5905_ _0736_ _0737_ _1070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_81_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6885_ _2009_ _0097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5648__I _0345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4552__I _3122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8624_ _0112_ clknet_4_0_0_Clock C\[0\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5836_ _0310_ _4137_ _1002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8555_ _0000_ clknet_4_2_0_Clock A\[0\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5767_ _0336_ _0937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5923__A3 _0647_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7506_ _2623_ _2629_ _2656_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4718_ _4030_ _4038_ _4039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8486_ _3673_ _3667_ _3686_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5698_ C\[2\]\[0\] _3870_ _4239_ _0462_ _0871_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_107_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4649_ _3854_ _3971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7437_ _2573_ _2582_ _2583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7676__A3 _2829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7368_ _2423_ _2426_ _2508_ _2509_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6319_ _0031_ _0054_ _1469_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7299_ _1018_ _2257_ _2434_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5439__A2 _0354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6939__A2 _2001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7061__A1 _2051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7364__A2 _2504_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6167__A3 _4093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8313__A1 _3461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5127__A1 _4033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6875__A1 _3798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7052__A1 _2049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5602__A2 _0203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4372__I _3229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6670_ _1722_ _1751_ _1799_ _1804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8552__A1 _0093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5621_ _0476_ _0795_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8340_ _3536_ _3538_ _3539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5552_ _0636_ _0640_ _0729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8304__A1 _3496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7107__A2 _1863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4503_ _3814_ _3818_ _3825_ _3826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5118__A1 _0178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8271_ _3463_ _3403_ _3464_ _3465_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5483_ C\[2\]\[7\] _3860_ _3928_ _0658_ _0660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_133_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5669__A2 C\[2\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6866__A1 _3949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7222_ _3817_ _2350_ _2351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4434_ _3752_ _3754_ _2341_ _3756_ _3757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_99_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6330__A3 _0469_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7153_ _3982_ C\[1\]\[8\] _2155_ _2275_ _2277_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4365_ _2971_ _3144_ _3163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6618__A1 _2816_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6104_ _0705_ _1263_ _1264_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6618__B2 A\[1\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7084_ _3889_ _2203_ _2125_ _2204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4296_ _2427_ _2438_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6035_ _1194_ _1197_ _1198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4547__I _3860_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7291__A1 _3968_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6094__A2 _0651_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xrebuffer10 _1713_ net43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_39_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7986_ _0049_ _0014_ _3071_ _3156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7594__A2 _2746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6937_ _2042_ _2059_ _2060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4282__I net4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6868_ _3957_ _1725_ _1992_ _1993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8543__A1 _0106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7346__A2 _1952_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8607_ _0052_ clknet_4_1_0_Clock B\[2\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5357__A1 _3842_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5819_ _0978_ _0979_ _0984_ _0985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5357__B2 _4169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6799_ A\[1\]\[5\] _1926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8538_ _0120_ _0075_ _0105_ _0090_ _3678_ _3719_ _3731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_109_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5109__A1 _0281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5327__B B\[0\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8469_ _3663_ _3667_ _3668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6857__A1 _3260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6321__A3 _1358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4332__A2 net7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4885__C _4200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6085__A2 _1099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7282__A1 _2400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6388__A3 _1534_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5288__I _0460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4406__B _3593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8534__A1 _0103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5348__A1 _0418_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4571__A2 net12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5520__A1 _0645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4323__A2 _2717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5751__I _0358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7273__A1 _3873_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4367__I _2330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7273__B2 _2053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5823__A2 _4188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7025__A1 _2085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7840_ _0344_ _1863_ _3001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7771_ _4158_ _0751_ _2237_ _2928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4983_ _4248_ _4249_ _4235_ _0169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_75_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6722_ _1836_ _1853_ _1854_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8525__A1 _3719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5339__A1 _0512_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6653_ _3402_ _1707_ _1787_ _1788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6000__A2 _3760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5604_ _3814_ _0383_ _0778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6584_ _1705_ _1720_ _1722_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8323_ _0457_ C\[0\]\[12\] _3521_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5535_ _3973_ C\[2\]\[9\] _0712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6839__A1 _3004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5466_ _0560_ _0580_ _0643_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8254_ _3442_ _3446_ _3447_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7205_ _2179_ _1757_ _2239_ _2333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4417_ _3701_ _3709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5511__A1 _0027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5397_ _3896_ _0574_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_82_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8185_ _0750_ _2013_ _2102_ _0051_ _3372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4348_ _2805_ net9 _2982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7136_ _3817_ _2257_ _2258_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4277__I net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7264__A1 _2334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7067_ _2178_ _2182_ _2187_ _2188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_4279_ _2244_ _2254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_87_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6018_ _3925_ _1181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4617__A3 _3938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8624__D _0112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5578__A1 _0201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7969_ _3054_ _3057_ _3139_ _3140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8618__CLK clknet_4_7_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8516__A1 _0129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7319__A2 _2455_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6058__A2 _0687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7255__A1 _2320_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4650__I _3971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xrebuffer1 _1790_ net34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
X_5320_ _0494_ _0495_ _0496_ _0497_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_6_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6577__I _1715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5251_ _3890_ net5 _0430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_47_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5182_ _0362_ _0363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_68_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_7_0_Clock_I clknet_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7797__A2 _2954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7823_ _2862_ _2981_ _2929_ _2927_ _2983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7754_ _2860_ _2865_ _2910_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4966_ _0149_ _0151_ _0152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6705_ _1247_ C\[1\]\[2\] _1723_ _1781_ _1837_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_51_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6261__B _1412_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7685_ _2837_ _0125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4897_ _4209_ _4211_ _4212_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4560__I _3877_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6636_ _1770_ _1771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7721__A2 _1999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5732__A1 _0847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4535__A2 _3856_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6567_ _2244_ _2265_ _2383_ _1706_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_69_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8306_ _3497_ _3502_ _3503_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5518_ _0622_ _0669_ _0694_ _0695_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6498_ _1624_ _1625_ _1641_ _1642_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8237_ _3356_ _3357_ _3428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8619__D _0068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5449_ _0554_ _0555_ _0626_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_117_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8168_ _3270_ _3329_ _3353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7237__A1 _1178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7119_ _2238_ _2239_ _2240_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_87_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8099_ _3277_ _3191_ _3263_ _3278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7788__A2 _0388_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4735__I _4014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output23_I net23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6212__A2 _1250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7960__A2 _3128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8590__CLK clknet_4_2_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4774__A2 _4091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4470__I _3792_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7712__A2 _2865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5723__A1 _4073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5487__B1 _0662_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6451__A2 _1533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4462__A1 B\[1\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4462__B2 _3784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6860__I _3931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4820_ _3872_ _3122_ _4137_ _3859_ _4138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8053__S _3228_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4765__A2 _3764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4751_ _4071_ _4072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_14_0_Clock_I clknet_3_7_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4380__I _3315_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4682_ _3949_ _4003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7470_ _2617_ _2618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7703__A2 _2778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6421_ _1475_ _1489_ _1567_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6352_ _1500_ _1501_ _1502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5190__A2 _0370_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5303_ _0479_ _0480_ _0481_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7467__A1 _1538_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6283_ _0045_ _1037_ _1434_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8022_ _3109_ _3117_ _3195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_103_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5234_ _0353_ _0415_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5165_ _0330_ _0346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_68_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5096_ _0263_ _0274_ _0279_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6442__A2 _1501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8195__A2 _3382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7806_ _0278_ _0291_ _2966_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_13_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5998_ _1017_ _1033_ _1161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7737_ _2893_ _0111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4949_ _0027_ _3240_ _4263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7668_ _0435_ _0003_ _2822_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5705__A1 _0848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6619_ _1754_ _1755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7599_ _2748_ _2751_ _2752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_4_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7458__A1 _2103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8186__A2 _3372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4747__A2 _4067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5944__A1 _1100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5172__A2 _0352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8110__A2 _1809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6855__I _1971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6672__A2 _1798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4683__A1 _4001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4683__B2 _3979_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4375__I _3260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6424__A2 C\[2\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6970_ _2060_ _2092_ _2093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4435__A1 _3709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5921_ _0707_ _1084_ _1085_ _1086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6590__I _1726_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8640_ _0096_ clknet_4_0_0_Clock C\[1\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5852_ _3934_ _1018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7924__A2 _1929_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4803_ _4043_ _4100_ _4121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5935__A1 _0342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8571_ _0016_ clknet_4_6_0_Clock A\[2\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5783_ _0950_ _0951_ _0952_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_72_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7522_ _2612_ _2616_ _2618_ _2673_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4734_ _4054_ _4048_ _4055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7453_ _2560_ _2564_ _2600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4665_ _3959_ _3963_ _3986_ _3987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_134_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6404_ _1508_ _1550_ _1551_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_128_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7384_ _2523_ _2525_ _2526_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4596_ _3917_ _3814_ _3918_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6335_ _4161_ _0039_ _1485_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6266_ _1296_ _1300_ _1417_ _1418_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8005_ _3094_ _3175_ _3176_ _3177_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5217_ _0397_ _0398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_15_0_Clock clknet_3_7_0_Clock clknet_4_15_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_83_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6197_ _1234_ _1350_ _1351_ _1352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4674__A1 _3800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5148_ _2610_ _2265_ _0330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_85_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4285__I net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5079_ _0237_ _0245_ _0262_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4426__A1 _3746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6966__A3 _2088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6714__B A\[0\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4977__A2 _0151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8632__D _0106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5926__A1 _1037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8340__A2 _3538_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4901__A2 _4213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6103__A1 _1038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7851__A1 _0479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6654__A2 _1710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7851__B2 _1734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4968__A2 _0153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5917__A1 _1077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5393__A2 _0569_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5754__I _0924_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4450_ _3772_ _3773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6342__B2 _1365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4381_ _3240_ _3326_ _3337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6120_ _1131_ _1192_ _1279_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8095__A1 _3194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6585__I B\[1\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6051_ _1065_ _1211_ _1212_ _1213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7842__A1 _3793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5002_ _0183_ _0187_ _0188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_112_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4319__B _2674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7070__A2 _2170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6953_ _3562_ _1848_ _2076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5904_ _1066_ _1067_ _1068_ _1069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6884_ _1934_ _2008_ _2009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8623_ _0111_ clknet_4_0_0_Clock C\[0\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5835_ _0982_ _0999_ _1000_ _1001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_22_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8554_ _0132_ clknet_4_14_0_Clock net23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5766_ _0919_ _0932_ _0936_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8651__CLK clknet_4_11_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7505_ _2653_ _2633_ _2654_ _2655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4717_ _3869_ _4037_ _4038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8485_ _0066_ _3681_ _3684_ _0064_ _3685_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_120_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5697_ _0753_ _0831_ _0870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8322__A2 _3469_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8040__I _3018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7436_ _2576_ _2581_ _2582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4648_ _3965_ _3969_ _3970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6333__A1 _1375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4344__B1 _2930_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7367_ _2424_ _2425_ _2508_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_122_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4579_ _3889_ _3900_ _3901_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8086__A1 _3184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6318_ _1466_ _1467_ _1468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_46_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7298_ _2361_ _2431_ _2432_ _2433_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7833__A1 _2926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8627__D _0115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6249_ _0985_ _1127_ _1193_ _1401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8010__A1 _0529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5574__I _0750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5127__A2 _0308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6875__A2 _1999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8077__A1 _3160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7824__A1 _0838_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8326__S _3523_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5063__A1 _4263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5602__A3 _0378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8674__CLK clknet_4_4_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8552__A2 _3681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5620_ _0342_ _0498_ _0793_ _0794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_34_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5551_ _0636_ _0640_ _0728_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8304__A2 _3500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4502_ _3820_ _3822_ _3824_ _3825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__5118__A2 _0300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8270_ _3398_ _3400_ _3464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5482_ C\[2\]\[7\] _4242_ _0658_ _3860_ _0659_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_144_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7221_ _2164_ _2350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4433_ _3755_ _3756_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_104_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7152_ _1902_ _2275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4364_ _2971_ _3144_ _3152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4341__A3 _2287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6618__A2 _1742_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6103_ _1038_ _0036_ _1263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_115_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4295_ _2308_ _2416_ _2427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7083_ _2126_ _2203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4629__A1 _3948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6034_ _0975_ _1195_ _1196_ _1197_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5841__A3 _1006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer11 _3572_ net44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
XTAP_2209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8240__A1 _3368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7985_ _3077_ _3136_ _3154_ _3155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5054__A1 _0192_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6936_ _2043_ _2058_ _2059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6867_ _4087_ _1990_ _1992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8543__A2 _3714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8606_ _0051_ clknet_4_1_0_Clock B\[2\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5818_ _4028_ _0982_ _0983_ _4129_ _0984_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_52_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5357__A2 _0413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6798_ _1925_ _0096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8537_ _3730_ _0144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5394__I _0509_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5749_ _0336_ _3790_ _0920_ _0921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_108_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8468_ net13 _3667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6857__A2 _1848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7419_ _1538_ _2562_ _2563_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8399_ _1673_ _3599_ _3600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4868__A1 _3793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8059__A1 _3194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4738__I A\[2\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5293__A1 _0463_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8697__CLK clknet_4_7_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7990__B1 _3098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8534__A2 _3666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5348__A2 _0425_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7273__A2 _1810_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7025__A2 _2088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8222__A1 _3390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5479__I _0576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7770_ _0896_ _1814_ _2927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5587__A2 _0761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4982_ _0162_ _0166_ _0167_ _0168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6721_ _1837_ _1845_ _1852_ _1853_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_60_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8525__A2 _0101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6652_ A\[0\]\[2\] _1787_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5603_ _2706_ _0493_ _0777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6583_ _1721_ _0066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8289__A1 _3427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8322_ _3466_ _3469_ _3519_ _3520_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5534_ _0710_ _0711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6839__A2 _1747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8253_ _0444_ _1930_ _3446_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5465_ _0573_ _0642_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_105_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7204_ _2328_ _2331_ _2332_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4416_ _3691_ _3701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5511__A2 _0687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8184_ _3284_ _3370_ _3371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5396_ _0567_ _0570_ _0572_ _0573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_67_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7135_ _2185_ _2257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4347_ _2889_ _2963_ _2971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7066_ _2183_ _2184_ _2186_ _2187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_4278_ net3 _2244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_87_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6017_ _4045_ _4067_ _4179_ _1179_ _1180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_86_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8213__A1 _0633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5027__A1 _0201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5578__A2 _0052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7968_ _3060_ _3138_ _3139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6775__A1 _3971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6919_ _1964_ _1968_ _2042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7899_ _2983_ _2984_ _3063_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__8640__D _0096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5852__I _3934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8452__A1 _3627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4608__A4 _3929_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8204__A1 _3311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6766__A1 _3767_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7191__A1 _2248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xrebuffer2 _1874_ net35 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5250_ _4159_ _0023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4378__I _3293_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5181_ _0344_ _0362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5009__A1 C\[3\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7822_ _1753_ _0317_ _1755_ _2981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_92_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7753_ _2849_ _2811_ _2907_ _2909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4965_ _0150_ _4219_ _0151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6704_ _1834_ _1792_ _1835_ _1836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_75_1384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7684_ _0954_ _0955_ _2837_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4896_ _3510_ _0029_ _4210_ _4211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_138_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6635_ _1724_ _1770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6566_ _3809_ _0040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4535__A3 _3857_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4997__B _0182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8305_ _3498_ _3501_ _3502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5517_ _0625_ _0668_ _0694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6497_ _1639_ _1640_ _1641_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8236_ _3425_ _3426_ _3427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5448_ _0559_ _0623_ _0624_ _0625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6288__A3 _4176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5496__A1 _0587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8167_ _3274_ _3328_ _3352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5379_ _4168_ _0392_ _0556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7118_ _4214_ _2164_ _2239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8098_ _0308_ _1758_ _3275_ _3276_ _3277_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__5248__A1 _0406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7049_ _2144_ _2147_ _2169_ _2170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_41_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6996__A1 _2043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7945__B1 _0566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output16_I net16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4751__I _4071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6920__A1 _1974_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5723__A2 _0032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6678__I _1810_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5582__I _0436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5487__A1 _3875_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5487__B2 _0468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6987__A1 _2025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5411__A1 _0214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5411__B2 _0437_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4661__I _3982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4750_ _3751_ _4071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4681_ _3823_ _4002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7703__A3 _2829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6420_ _1477_ _1565_ _1566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6351_ _1394_ _1396_ _1392_ _1501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6588__I _1725_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5302_ _3456_ _3260_ _0350_ _0480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_143_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7467__A2 _2614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6282_ _1318_ _1327_ _1432_ _1433_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_1407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8021_ _3177_ _3179_ _3193_ _3194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_115_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5233_ _0413_ _0414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8608__CLK clknet_4_11_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7219__A2 _2261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5164_ _0344_ _0345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5095_ _0256_ _0276_ _0277_ _0278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7805_ _2965_ _0112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5997_ _1143_ _1159_ _1160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5402__A1 C\[2\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7736_ _2839_ _2892_ _2893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4948_ _4262_ _0027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5953__A2 _0747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_11_0_Clock clknet_3_5_0_Clock clknet_4_11_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_127_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7667_ _0924_ _1975_ _2821_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7155__A1 _1018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4879_ _4195_ _0059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6618_ _2816_ _1742_ _1743_ A\[1\]\[2\] _1754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_7598_ _2749_ _2750_ _2751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6549_ C\[3\]\[16\] _1628_ _1687_ _1690_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7458__A2 _2570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7831__B _2958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8219_ _3407_ _3408_ _3409_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_106_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6130__A2 _1189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6969__A1 _2064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7394__A1 _2411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4747__A3 _3950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7146__A1 _4001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7697__A2 _2811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7449__A2 _2581_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6121__A2 _1192_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4656__I _3812_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4683__A2 _3778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6424__A3 B\[2\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5632__A1 _0804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4435__A2 _3751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5920_ _0709_ _0723_ _1085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5851_ _4175_ _4186_ _1016_ _1017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4802_ _4109_ _4119_ _4120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_34_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8570_ _0015_ clknet_4_3_0_Clock A\[1\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5782_ _0016_ _0757_ _0951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5935__A2 _1099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7521_ _2658_ _2671_ _2672_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4733_ _3825_ _3951_ _4054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7137__A1 _3968_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7452_ _2569_ _2583_ _2597_ _2598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4664_ _3970_ _3977_ _3985_ _3986_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6403_ _1509_ _1549_ _1550_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7383_ _2456_ _2463_ _2525_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4595_ _3916_ _3917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6334_ _1483_ _1484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6265_ _0061_ _3646_ _1301_ _1417_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_142_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8004_ _3090_ _3097_ _3176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_83_1461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5216_ _3840_ _0397_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6196_ _0054_ _1234_ _1351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4674__A2 _0042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8580__CLK clknet_4_1_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5147_ _0324_ _0328_ _0329_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_111_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6415__A3 _1358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7612__A2 _1704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5078_ _0237_ _0245_ _0261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input15_I reset vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4426__A2 _3748_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6820__B1 _1761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6179__A2 _1335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5397__I _3896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4515__B A\[3\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5926__A2 _0403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4729__A3 _3986_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7719_ _0922_ _0923_ _1847_ _1850_ _4066_ _2874_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__7128__A1 _4076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8699_ _0145_ clknet_4_13_0_Clock net19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6887__B1 _1698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6021__I _3992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4901__A3 _4215_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7300__A1 _0473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6103__A2 _0036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7851__A2 _0480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5862__A1 _3777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4665__A2 _3963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4476__I _3798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4380_ _3315_ _3326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6050_ _1069_ _1113_ _1212_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_113_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7842__A2 _0751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input7_I X[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4386__I _3380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5853__A1 _3761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5001_ C\[3\]\[1\] _0186_ _0187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6952_ _2745_ _1777_ A\[0\]\[6\] _2075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5903_ _0698_ _0724_ _1068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6883_ _1937_ _2007_ _2008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__7358__A1 _4090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5834_ _3849_ _3615_ _1000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8622_ _0110_ clknet_4_1_0_Clock C\[0\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5765_ _0919_ _0932_ _0935_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8553_ _3645_ _3687_ _3742_ _3743_ _0148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_124_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6581__A2 _1718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4716_ _3868_ _4032_ _4036_ _4037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_7504_ _2611_ _2632_ _2654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8484_ _3683_ _3674_ _3684_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5696_ _0868_ _0869_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5166__B B\[0\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7435_ _2577_ _2580_ _2581_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_11_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4647_ _3968_ _3969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6333__A2 _1482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4344__A1 _2897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7366_ _2495_ _2506_ _2507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4578_ _3899_ _3900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8477__B _3671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6317_ _1354_ _1386_ _1467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7297_ _2364_ _2368_ _2432_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6248_ _1199_ _1202_ _1336_ _1399_ _1400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__8491__C1 _3676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7833__A2 _2931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5844__A1 _0998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6179_ _1281_ _1335_ _1336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_58_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7597__A1 _0048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8643__D _0099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8010__A2 _1928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4335__A1 _2794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8077__A2 _3166_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5590__I _0423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6088__A1 _3842_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7824__A2 _1952_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5835__A1 _0982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5602__A4 _0775_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4810__A2 _3844_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5550_ _0611_ _0619_ _0726_ _0727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4501_ _3823_ _3824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5481_ _0657_ _0658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7220_ _4035_ _1757_ _2349_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4432_ _3727_ _2373_ _2394_ _3755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_126_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6866__A3 _1990_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6596__I _1707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7151_ _2162_ _2165_ _2273_ _2274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4363_ _3026_ _3133_ _3144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6079__A1 _1098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6102_ _1260_ _1107_ _1261_ _1262_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7082_ _4116_ _0014_ _2122_ _2202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4294_ _2341_ _2405_ _2416_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4629__A2 _3937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6033_ _0977_ _1045_ _1196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7579__A1 _1597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer12 _0311_ net45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8240__A2 _3384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7984_ _3081_ _3135_ _3154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6935_ _2044_ _2049_ _2057_ _2058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_70_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6866_ _3949_ _1724_ _1990_ _1991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_126_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8605_ _0050_ clknet_4_0_0_Clock B\[2\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5817_ _4128_ _4131_ _0983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6797_ _1871_ _1872_ _1924_ _1925_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_50_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4565__A1 _3837_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8536_ _0119_ _0074_ _0104_ _0089_ _3678_ _3719_ _3730_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5748_ _0334_ _0920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8467_ _3665_ _3666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5679_ _0850_ _0851_ _0852_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7418_ _2163_ _2562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8398_ _1597_ C\[0\]\[14\] _3599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4868__A2 _3937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8059__A2 _3198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8638__D _0087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7349_ _2410_ _2487_ _2488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6490__A1 _1481_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7990__A1 _3000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5596__A3 _0361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4703__B _4017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7742__A1 _2842_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5808__A1 _0031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6481__A1 _1561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8641__CLK clknet_4_0_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4981_ _0163_ _0164_ _0165_ _0167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7981__A1 _3066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6720_ _4012_ _1851_ _1852_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_36_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6651_ _1782_ _1785_ _1786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5602_ _0774_ _0203_ _0378_ _0775_ _0776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_108_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6582_ _1705_ _1720_ _1721_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8321_ _3518_ _0005_ _3470_ _3519_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5533_ _0656_ _0710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8252_ _3290_ _3442_ _3443_ _3444_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5464_ _0629_ _0636_ _0640_ _0641_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_7203_ _2313_ _2329_ _2331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4415_ _2481_ net15 _3691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4839__I _4009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8183_ _0750_ _2101_ _3370_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5395_ _3953_ _0571_ _0572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7134_ _2253_ _2153_ _2255_ _2256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4346_ _2952_ _2963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7065_ _4214_ _2185_ _2186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4277_ net1 _2233_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__8461__A2 _0181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6472__A1 _1590_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6016_ _1178_ C\[3\]\[10\] _1179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8213__A2 _2250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5027__A2 _0211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6224__A1 _1037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7967_ _3062_ _3137_ _3138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5578__A3 _0753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6775__A2 C\[1\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4786__A1 _3902_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6918_ _1970_ _2004_ _2040_ _2041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7898_ _2989_ _3040_ _3061_ _3062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_1065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7724__A1 _0035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6849_ _1839_ _1975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4538__A1 _3260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4538__B2 B\[3\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8519_ _0099_ _3693_ _3713_ _3714_ _3715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_87_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4749__I _3955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8664__CLK clknet_4_15_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6964__I _2086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6215__A1 _0981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7963__A1 _3103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6766__A2 _1894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4777__A1 _3961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7191__A2 _2286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer3 _1821_ net36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_5_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4659__I _3980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5180_ _4072_ _0360_ _0361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6874__I _1998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6454__A1 _1598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5009__A2 _0184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6206__A1 _1245_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7821_ _2925_ _2932_ _2980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_58_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7954__A1 _0389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7752_ _2761_ _0012_ _2850_ _2907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4964_ _3791_ _4220_ _4216_ _3774_ _0150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6703_ _1833_ _1782_ _1785_ _1835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_51_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7683_ _2835_ _0080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4895_ _4206_ _4208_ _4210_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7706__A1 _2819_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6634_ _1768_ _1702_ _1769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6565_ _0208_ _1704_ _1705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5732__A3 _0873_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8304_ _3496_ _3500_ _3501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8687__CLK clknet_4_5_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5516_ _0682_ _0692_ _0693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_121_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6496_ _1626_ _1627_ _1638_ _1640_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__8131__A1 _1672_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5447_ _0563_ _0581_ _0624_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8235_ _3351_ _3418_ _3426_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8166_ _3349_ _3350_ _3351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5378_ _3751_ _0400_ _0555_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_59_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4329_ _2556_ _2786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7117_ _2236_ _2179_ _2237_ _2238_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_82_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8097_ _2998_ _3186_ _3276_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7048_ _2154_ _2158_ _2168_ _2169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_86_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6996__A2 _2058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8198__A1 _3366_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7945__A1 _3434_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7945__B2 _1770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8651__D _0093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5184__A1 _0356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6920__A2 _1976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8122__A1 _0392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5487__A2 _0658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6684__A1 _1815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6694__I _1826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6436__A1 _1561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6987__A2 _2094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8189__A1 _3189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7936__A1 _2871_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8561__D _0006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5411__A2 _0327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4680_ _3820_ _4001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_119_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8361__A1 _3518_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6911__A2 _1952_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6350_ _1388_ _1391_ _1500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4922__A1 _4222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8113__A1 _3286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5301_ _3531_ _2786_ _0330_ B\[0\]\[5\] _0479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_142_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4389__I _3413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6281_ _1321_ _1430_ _1431_ _1432_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_66_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5478__A2 _0654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6675__A1 _3776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8020_ _3184_ _3192_ _3193_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5232_ _0362_ _0413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5163_ _0343_ _0344_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8416__A2 _3541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6427__A1 _1481_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5094_ _0259_ _0275_ _0277_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4338__B _2867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5013__I _3133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7927__A1 _3091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7804_ _2898_ _2901_ _2964_ _2965_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_91_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5996_ _1145_ _1158_ _1159_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5402__A2 _4242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7735_ _2842_ _2891_ _2892_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4947_ _3845_ _4262_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7666_ _0823_ _1783_ _2820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4878_ _2963_ _4195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7155__A2 _2275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5166__A1 _2492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6617_ _2867_ _1753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7597_ _0048_ _0009_ _2750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4913__A1 _4227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6548_ _1688_ C\[3\]\[16\] _1689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8104__A1 _0314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4299__I net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6479_ _1623_ _0077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6666__A1 _1738_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8218_ _0488_ _3302_ _3408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8646__D _0088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8149_ _3060_ _3138_ _3333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_59_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6969__A2 _2091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7091__A1 _3004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8702__CLK clknet_4_13_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5641__A2 _0787_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7394__A2 _2473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7146__A2 _1319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4904__A1 _4218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6657__A1 _0179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8556__D _0001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7082__A1 _4116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6424__A4 _3898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4435__A3 _3757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7909__A1 _2760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5850_ _4178_ _1014_ _1015_ _1016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_62_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4801_ _4111_ _4115_ _4118_ _4119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_2190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5396__A1 _0567_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5781_ _0872_ _0949_ _0950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7520_ _2661_ _2670_ _2671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_72_1366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4732_ _4051_ _4016_ _4052_ _4053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7137__A2 _1841_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8334__A1 _3495_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7451_ _2548_ _2568_ _2597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4663_ _3979_ _3981_ _3984_ _3985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_119_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6402_ _1511_ _1548_ _1549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6896__A1 _1939_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7382_ _2452_ _2455_ _2523_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4594_ _3915_ _3753_ _3802_ _3755_ _3916_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6333_ _1375_ _1482_ _1483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_143_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6264_ _1414_ _1415_ _1416_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5215_ _0385_ _0394_ _0395_ _0396_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8003_ _3090_ _3097_ _3175_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6195_ _0030_ _0054_ _1350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7223__I _1962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5146_ _0206_ _0326_ _0328_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4674__A3 _3806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5077_ _0251_ _0260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7612__A3 _0010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6820__A1 _4202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6820__B2 _4195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5979_ _1001_ _1008_ _1142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7718_ _0348_ _0352_ _2871_ _2872_ _2236_ _2873_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_139_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8698_ _0144_ clknet_4_12_0_Clock net18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7128__A2 _0004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5139__A1 _3875_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7649_ _2799_ _2800_ _2801_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6887__A1 _2010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6887__B2 _3967_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_9_0_Clock clknet_3_4_0_Clock clknet_4_9_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_101_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7300__A2 C\[1\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4757__I _3787_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5862__A2 _3789_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4665__A3 _3986_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5614__A2 _0787_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6811__A1 _1815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4492__I B\[1\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5378__A1 _3751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8316__A1 _3465_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6878__A1 _1974_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5302__A1 _3456_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7043__I _2163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7842__A3 _3002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5000_ _0185_ _0186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5853__A2 _4168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7055__A1 _2438_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5066__B1 _0220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6951_ _1985_ _1894_ _2074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5902_ _0744_ _1067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6882_ _1939_ _1942_ _2006_ _2007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_50_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7358__A2 C\[1\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8621_ _0102_ clknet_4_1_0_Clock C\[0\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5833_ _2460_ _3897_ _0999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6030__A2 _1192_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8552_ _0093_ _3681_ _3743_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5764_ _0916_ _0919_ _0932_ _0933_ _0934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_124_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7503_ _2607_ _2653_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4715_ _4033_ _4035_ _4036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8483_ _3663_ _3683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5695_ _0020_ _0757_ _0868_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7434_ _0062_ _2579_ _2402_ _2580_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4646_ _3966_ _3764_ _3967_ _3765_ _3968_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_129_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4344__A2 _2919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4577_ _3898_ _3899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7365_ _2500_ _2505_ _2506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8477__C _3676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6316_ _1356_ _1465_ _1466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7296_ _2364_ _2368_ _2431_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4577__I _3898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7294__A1 _2359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6247_ _1194_ _1197_ _1399_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8491__B1 _3684_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8491__C2 _0067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6178_ _1282_ _1334_ _1335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7046__A1 _2160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5129_ _0303_ _0311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_57_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7597__A2 _0009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7349__A2 _2487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8512__I _3686_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5780__A1 _0946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5532__A1 _0655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4335__A2 _2826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5871__I _4062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7760__A2 _2915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5771__A1 _0928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8570__CLK clknet_4_3_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4500_ A\[2\]\[1\] _3787_ _3797_ _3788_ _3823_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_5480_ _0656_ _0657_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4431_ _3753_ _3754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5523__A1 _0637_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4362_ _3122_ _3133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7150_ _4090_ C\[1\]\[7\] _2156_ _1840_ _2273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_98_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7276__A1 _2403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6101_ _1105_ _1106_ _1261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_112_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7081_ _2130_ _2199_ _2200_ _2201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4293_ _2352_ _2373_ _2394_ _2405_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_98_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4629__A3 _3950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6032_ _0977_ _1045_ _1195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7028__A1 _1985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7579__A2 C\[0\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7983_ _3150_ _3151_ _3153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6934_ _2051_ _2052_ _2056_ _2057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__5021__I _4033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6865_ _3982_ C\[1\]\[5\] _1990_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7200__A1 _2252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6003__A2 _1023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8604_ _0049_ clknet_4_1_0_Clock B\[2\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5816_ _0980_ _0981_ _0982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6796_ _1815_ _1874_ _1923_ _1924_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_8535_ _3726_ _3728_ _3729_ _0143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5747_ _0910_ _0911_ _0895_ _0919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__5762__A1 _0921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8466_ _3663_ _3664_ _3665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5678_ _0791_ _0798_ _0851_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_136_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5514__A1 _0689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4317__A2 _2652_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7417_ _1295_ _1930_ _2561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4629_ _3948_ _3937_ _3950_ _3951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_8397_ _3556_ _3558_ _3597_ _3598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4868__A3 _3980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7348_ _2484_ _2486_ _2487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_137_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7279_ _0060_ _2013_ _2102_ _0059_ _2412_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7019__A1 _3816_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8519__A1 _0099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8593__CLK clknet_4_10_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4770__I _4089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4556__A2 _3878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5505__A1 _0589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_3_6_0_Clock clknet_0_Clock clknet_3_6_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_122_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5808__A2 _0057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8564__D _0009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4980_ _0163_ _0164_ _0165_ _0166_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_45_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7981__A2 _3075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6784__A3 _1912_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4680__I _3820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6650_ _4157_ _1783_ _1784_ _1785_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_31_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5601_ _0389_ _0775_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5744__A1 _0914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6581_ _1717_ _1718_ _1719_ _1720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8320_ _0506_ _3518_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5532_ _0655_ _0666_ _0708_ _0709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8251_ _0053_ _1931_ _3379_ _3443_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5463_ _0637_ _0638_ _0639_ _0640_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_7202_ _4195_ _2012_ _2329_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4414_ _3347_ _3672_ _3682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8182_ _3204_ _3205_ _3323_ _3367_ _3368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_99_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5394_ _0509_ _0571_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_114_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7133_ _2148_ _2149_ _2255_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_119_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4345_ _2941_ _2952_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5016__I _0201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7064_ _2086_ _2185_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6015_ _3890_ _1178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4855__I _4172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6224__A2 _0037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7966_ _3077_ _3136_ _3137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6917_ _1973_ _2003_ _2040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5983__A1 _3844_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7897_ _2992_ _3039_ _3061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6848_ _1896_ _1900_ _1974_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_52_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7724__A2 _1716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5735__A1 _0848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4538__A2 _2919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6779_ _3767_ _1907_ _1904_ _0476_ _1908_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_109_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8518_ _3665_ _3714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7488__A1 _2544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8649__D _0091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8449_ C\[0\]\[16\] _1628_ _3651_ _3653_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_100_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6160__A1 _0044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7660__A1 _2811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6215__A2 _0711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6980__I _2101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7412__A1 _2552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6766__A3 _1842_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4777__A2 _3824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrebuffer4 net41 net37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_122_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8559__D _0004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6890__I _2013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7820_ _2916_ _2917_ _2978_ _2979_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7954__A2 _1962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7751_ _2854_ _2888_ _2905_ _2906_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4963_ _4272_ _4274_ _4276_ _0149_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_36_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6702_ _1782_ _1785_ _1833_ _1834_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7682_ _0228_ _0254_ _2835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4894_ _4206_ _4208_ _4209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7706__A2 _2823_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6633_ _2427_ _1768_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6564_ _1703_ _1704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8303_ _0445_ _2579_ _3500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5515_ _0684_ _0691_ _0692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6495_ _1626_ _1627_ _1638_ _1639_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8131__A2 _3312_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8234_ _3354_ _3417_ _3425_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5446_ _0563_ _0581_ _0623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8165_ _3262_ _3269_ _3350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5377_ _3604_ _0376_ _0554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_99_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7116_ _1754_ _2237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4328_ _2745_ _2755_ _2764_ A\[3\]\[2\] _2775_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_99_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8096_ _3088_ _3096_ _3275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7047_ _2166_ _2167_ _2168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5956__A1 _0866_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7949_ _3023_ _3109_ _3117_ _3118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8370__A2 _0014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8631__CLK clknet_4_10_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5184__A2 _3848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8122__A2 _3302_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4695__A1 _4012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4495__I _3817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8189__A2 _3375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7936__A2 _2872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7164__A3 _2288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8361__A2 _2665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6372__A1 _1300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8113__A2 _3289_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5300_ _0475_ _0477_ _0478_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6280_ _1323_ _1324_ _1326_ _1431_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5231_ _0407_ _0410_ _0411_ _0412_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_45_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7872__A1 _3028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6885__I _2009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6675__A2 _1807_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5162_ _2816_ _0311_ _0312_ B\[2\]\[2\] _0343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__7624__A1 _2772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5093_ _0259_ _0275_ _0276_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7927__A2 _3093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7803_ _2904_ _2962_ _2964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_52_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5938__A1 _0800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5995_ _1157_ _1158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5938__B2 _3976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8541__S _3695_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7734_ _2799_ _2846_ _2890_ _2891_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_4946_ _4194_ _4260_ _4261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8654__CLK clknet_4_4_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4610__A1 _3931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7665_ _2817_ _2776_ _2818_ _2819_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_1284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4877_ _3911_ _4193_ _4194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_127_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6616_ _1752_ _0067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5166__A2 _3782_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7596_ _0375_ _1704_ _2749_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_14_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6547_ _1598_ _1688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4913__A2 _3905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8104__A2 _2011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6478_ _1617_ _1622_ _1623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_84_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8217_ _0720_ _1987_ _3407_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5429_ _0552_ _0558_ _0605_ _0606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8148_ _3253_ _3331_ _3332_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_59_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7615__A1 _2733_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6418__A2 _1492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8079_ _3158_ _3254_ _3255_ _3256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_87_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7091__A2 _1814_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8662__D _0131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_5_0_Clock clknet_3_2_0_Clock clknet_4_5_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_43_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7146__A3 _1980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8343__A2 _3541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4904__A2 _3809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7854__A1 _3013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6657__A2 _1791_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7606__A1 _0375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7082__A2 _0014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8677__CLK clknet_4_12_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7909__A2 _2203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8031__A1 _0924_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4800_ _4107_ _4117_ _4118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5780_ _0946_ _0948_ _0949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6593__A1 _1727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4731_ _4008_ _4011_ _4052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_30_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7450_ _2573_ _2582_ _2595_ _2596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4662_ _3983_ C\[3\]\[6\] _3984_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5148__A2 _2265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6401_ _1522_ _1547_ _1548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7381_ _2466_ _2521_ _2522_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_134_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4593_ B\[1\]\[4\] _3915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8098__A1 _0308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6332_ _1478_ _1480_ _1481_ _1482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7845__A1 _2997_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6263_ _0060_ _3900_ _1303_ _1415_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8002_ _3103_ _3171_ _3172_ _3134_ _3099_ _3173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_131_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5214_ _4275_ _0374_ _0377_ _0384_ _0395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5320__A2 _0495_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6194_ _0687_ _0054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5145_ _0326_ _0327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5076_ _0210_ _0257_ _0258_ _0259_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6820__A2 _1740_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8022__A1 _3109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5387__A2 _2578_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5978_ _1004_ _1007_ _1141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7781__B1 _1847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7717_ _2826_ _1848_ _2872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4929_ _3918_ _3923_ _4243_ _4244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_8697_ _0143_ clknet_4_7_0_Clock net17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8325__A2 _2087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7648_ _2761_ _1748_ _1812_ _2797_ _2800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__6336__A1 _1038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6887__A2 _3776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7579_ _1597_ C\[0\]\[0\] _0757_ _0000_ _2733_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_119_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8657__D _0126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7836__A1 _2938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6639__A2 _1773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7836__B2 _2937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5862__A3 _4182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4773__I _4092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4822__A1 _2685_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8013__A1 _3947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5378__A2 _0400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6878__A2 _1976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8567__D _0012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5302__A2 _3260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5853__A3 _1018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7055__A2 _1927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5066__A1 _0027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5066__B2 _0026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5605__A3 _0394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6950_ _1989_ _2001_ _2072_ _2073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_19_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4813__A1 _3849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5901_ _0698_ _0724_ _1066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6881_ _1956_ _1959_ _2005_ _2006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_78_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7358__A3 _2156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8620_ _0069_ clknet_4_1_0_Clock C\[0\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5832_ _4153_ _4164_ _0997_ _0998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8551_ _3704_ _0123_ _3686_ _3741_ _3742_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5763_ _0914_ _0915_ _0933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7502_ _2603_ _2604_ _2605_ _2602_ _2651_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_4714_ _4034_ _4035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8482_ _3675_ _3681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5694_ _0857_ _0859_ _0867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_0_Clock Clock clknet_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_124_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6869__A2 _1993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7433_ _2123_ _2579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4645_ _3413_ net11 _3967_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7364_ _2502_ _2504_ _2505_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4576_ _3897_ _3898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6315_ _1359_ _1385_ _1465_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7295_ _2422_ _2429_ _2430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6246_ _1398_ _0120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8491__A1 _0069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7294__A2 _2428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8491__B2 _0065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6177_ _1284_ _1333_ _1334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_97_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5128_ _4031_ _0310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8243__A1 _3371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5057__A1 _0193_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4593__I B\[1\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5059_ _4113_ _0200_ _0242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4335__A3 _2836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4768__I _4087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6088__A3 _1248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5296__A1 _0473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8234__A1 _3354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7037__A2 _2088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6796__A1 _1815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6548__A1 _1688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_2_0_Clock clknet_0_Clock clknet_3_2_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_44_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4430_ _2737_ _3746_ _3747_ _2567_ _3753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_144_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6720__A1 _4012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5523__A2 _0638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6379__B _1438_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4678__I _3998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4361_ _3111_ _3122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_67_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6100_ _1105_ _1106_ _1260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_125_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7080_ _2132_ _2191_ _2200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7276__A2 _2408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4292_ _2383_ _2394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_119_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5287__A1 _0398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6031_ _1128_ _1193_ _1194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7028__A2 _1907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7579__A3 _0757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7982_ _3064_ _3076_ _3151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6933_ _2053_ _2055_ _2056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6864_ _1984_ _1988_ _1989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5815_ _3315_ _0981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8603_ _0048_ clknet_4_0_0_Clock B\[2\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6795_ _1877_ _1913_ _1922_ _1923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_50_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8534_ _0103_ _3666_ _3729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5746_ _0888_ _0916_ _0917_ _0918_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8465_ net13 _3664_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5677_ _0841_ _0846_ _0849_ _0850_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7416_ _2502_ _2560_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4628_ _3949_ _3950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6711__A1 _1838_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8396_ _3518_ _0007_ _3559_ _3597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7347_ _3877_ _2120_ _2485_ _2486_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4559_ _3870_ _3882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7278_ _2329_ _2410_ _2411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6229_ _1379_ _1380_ _1381_ _1382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_131_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8216__A1 _0390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5212__I _0392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5450__A1 _4080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8519__A2 _3693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8670__D _0064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8523__I _3717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6950__A1 _1989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6978__I _2099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4498__I _2867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4713__B1 _3893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7258__A2 _2340_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8207__A1 _3312_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6769__A1 _3819_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5122__I _0303_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5441__A1 _0615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8580__D _0025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4961__I _3965_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5992__A2 _1153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7718__B1 _2871_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5600_ _3964_ _0774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6580_ _1479_ C\[1\]\[0\] _0040_ _1715_ _1719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__6941__A1 _1979_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6941__B2 _2043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5531_ _0661_ _0665_ _0708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6888__I _2011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8250_ _1099_ _1949_ _3442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7497__A2 _2646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5462_ _0422_ _0393_ _0639_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7201_ _1768_ _2100_ _2328_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4413_ _0056_ _0030_ _3662_ _3672_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8181_ _0899_ _2614_ _3367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5393_ _3921_ _0569_ _0570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7132_ _2148_ _2149_ _2253_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4344_ _2897_ _2919_ _2930_ B\[3\]\[3\] _2941_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_67_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7063_ _3821_ _3866_ _2050_ _2184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_80_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6014_ _1029_ _1031_ _1176_ _1177_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7965_ _3081_ _3135_ _3136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_36_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5432__A1 _4130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6916_ _2028_ _2038_ _2039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_70_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5983__A2 _0574_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7896_ _3058_ _3059_ _3060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6847_ _3962_ _1972_ _1911_ _1910_ _1893_ _1973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__7185__A1 _2223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7724__A3 _2824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6778_ _1903_ _1907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6798__I _1925_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8517_ _3692_ _3711_ _3712_ _3713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5729_ _0898_ _0900_ _0825_ _0901_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_143_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8448_ _1688_ C\[0\]\[16\] _3652_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_108_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8379_ _3495_ _3548_ _3578_ _3533_ _3493_ _3579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_102_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6160__A2 _4062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8665__D _0120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5671__A1 _0342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8560__CLK clknet_4_10_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5423__A1 _0548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4777__A3 _4096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6923__A1 _4112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5726__A2 _0897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer5 _1780_ net38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8575__D _0020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6454__A3 _1534_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5662__A1 _0833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4465__A2 _3445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7403__A2 _2506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4691__I _3832_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7750_ _2858_ _2887_ _2905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4962_ _4275_ _4215_ _4220_ _4276_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5965__A2 _1044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6701_ _1374_ C\[1\]\[1\] _1723_ _0000_ _1833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7681_ _2834_ _0110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4893_ _0028_ _3240_ _4208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6632_ _1760_ _1764_ _1766_ _1767_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_6563_ _1702_ _1703_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5514_ _0689_ _0690_ _0691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8302_ _0053_ _2203_ _3498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6494_ _1632_ _1634_ _1637_ _1638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_8233_ _3343_ _3420_ _3422_ _3424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_69_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5445_ _0604_ _0621_ _0622_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6142__A2 _1300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8164_ _3266_ _3268_ _3349_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5376_ _0507_ _0510_ _0553_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7115_ _1753_ _2236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5471__B _3946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8583__CLK clknet_4_4_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4327_ _2524_ _2764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_141_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8095_ _3194_ _3272_ _3273_ _3274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7046_ _2160_ _2162_ _2165_ _2167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5653__A1 _4275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7945__A3 _1181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8073__I _3238_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7948_ _3018_ _3115_ _3116_ _3117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_43_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5956__A2 _0964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7879_ _2901_ _2964_ _3044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5708__A2 _0880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5184__A3 _0364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_1_0_Clock clknet_3_0_0_Clock clknet_4_1_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_139_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4695__A2 _4015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4776__I _3980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7152__I _1902_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5400__I _0576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5230_ _2717_ _0315_ _0411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_29_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4686__I _3757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5161_ _0310_ _0342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_38_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5092_ _0248_ _0263_ _0274_ _0275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__7997__I _3022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7388__A1 _2457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7802_ _2906_ _2961_ _2962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5399__B1 _0306_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5994_ _1149_ _1156_ _1157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5310__I _0487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4945_ _4232_ _4258_ _4259_ _4260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7733_ _2854_ _2888_ _2890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4610__A2 _3761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4876_ _4105_ _4192_ _4193_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7664_ _2815_ _2773_ _1771_ _1972_ _2818_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_60_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6615_ _1722_ _1751_ _1752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7595_ _2733_ _2747_ _2748_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5166__A3 _0346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4374__A1 _2805_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6546_ C\[3\]\[15\] _1596_ _1599_ _1687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6477_ _1619_ _1621_ _1622_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6115__A2 _1119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8216_ _0390_ _2152_ _3406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5428_ _0507_ _0510_ _0557_ _0605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5874__A1 _0042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8147_ _3257_ _3261_ _3330_ _3331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_102_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5359_ _0534_ _0424_ _0535_ _0536_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8078_ _3160_ _3166_ _3255_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_59_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7029_ _3854_ _1777_ A\[0\]\[7\] _2150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7091__A3 _2208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5220__I _0400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4601__A2 _3922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7146__A4 _1999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7147__I _2269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4365__A1 _2971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6986__I _2022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7303__A1 _2367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6106__A2 _1265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7854__A2 _3014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5865__A1 _4045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7606__A2 _1748_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5617__A1 _0776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7610__I _2760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6290__A1 _0335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8031__A2 _2404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5130__I _0305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7790__A1 C\[0\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6593__A2 _1729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4730_ _4008_ _4011_ _4051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4661_ _3982_ _3983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6400_ _1543_ _1546_ _1547_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_70_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7380_ _2467_ _2469_ _2520_ _2521_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_4592_ _3811_ _3835_ _3914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_128_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6331_ _1374_ C\[2\]\[13\] B\[2\]\[7\] _3625_ _1481_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_128_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8098__A2 _1758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6262_ _1298_ _1302_ _1414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7845__A2 _3006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5856__A1 _1019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8001_ _3118_ _3132_ _3172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5213_ _0386_ _0393_ _0394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6193_ _1347_ _1348_ _1349_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5144_ _0325_ _0326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5608__A1 _0366_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5075_ _0234_ _0252_ _0258_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8621__CLK clknet_4_1_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5977_ _1011_ _1043_ _1139_ _1140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7781__A1 _0348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5387__A3 _0346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6584__A2 _1720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7781__B2 _1850_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7716_ _3037_ _1731_ A\[0\]\[2\] _2871_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_100_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4928_ C\[3\]\[4\] _4242_ _4243_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8696_ _0142_ clknet_4_13_0_Clock net32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7647_ _2760_ _1762_ _1814_ _2797_ _2799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_4859_ _4092_ _4176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6336__A2 _0038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4347__A1 _2889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7578_ _0048_ _0008_ _2732_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6529_ C\[2\]\[16\] _1671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8089__A2 _1928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5847__A1 _4165_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5862__A4 _1027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8673__D _0080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4822__A2 _3862_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8013__A2 _0576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6327__A2 _1376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4338__A1 _2775_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4889__A2 _4204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5838__A1 _3868_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8644__CLK clknet_4_8_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4510__A1 _3831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8583__D _0028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6263__A1 _0060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5066__A2 _0056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4813__A2 _4130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5900_ _0689_ _1064_ _1065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_34_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6880_ _1970_ _2004_ _2005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7358__A4 _2164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5831_ _4156_ _4163_ _0997_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_61_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8550_ _1666_ _1667_ _3675_ _3670_ _3741_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5762_ _0921_ _0930_ _0931_ _0932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_50_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7501_ _2649_ _2639_ _2650_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4713_ B\[3\]\[7\] _2930_ _3893_ _2919_ _4034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5693_ _0864_ _0865_ _0866_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8481_ _3660_ _3666_ _3677_ _3680_ _0132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7515__A1 _1597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4644_ B\[1\]\[6\] _3966_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7432_ _3883_ _2126_ _2577_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4575_ _3896_ _3897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7363_ _1319_ _1999_ _2152_ _1164_ _2504_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7279__B1 _2102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6314_ _1221_ _1462_ _1463_ _1464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7294_ _2359_ _2428_ _2429_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6245_ _1392_ _1397_ _1398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_143_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8491__A2 _3687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6176_ _1288_ _1291_ _1332_ _1333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_58_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5127_ _4033_ _0308_ _0309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5058_ _0239_ _0240_ _0195_ _0241_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA_input13_I Z[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6006__A1 _1028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8679_ _0086_ clknet_4_7_0_Clock C\[3\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7853__C _1753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8668__D _0123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8667__CLK clknet_4_15_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4740__B2 _3770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5296__A2 C\[2\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7745__A1 _2846_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5771__A3 _0921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8170__A1 _3281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8578__D _0023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4959__I _3953_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6720__A2 _1851_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4360_ _3056_ _3089_ _3100_ _3111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_125_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4291_ net4 _2383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_63_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6030_ _1131_ _1192_ _1193_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5287__A2 _0461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I X[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4694__I _4014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5039__A2 _0221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7579__A4 _0000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7981_ _3066_ _3075_ _3150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7984__A1 _3081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6932_ _2054_ _2055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6863_ _1985_ _1783_ _1987_ _4012_ _1988_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_63_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7736__A1 _2839_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8602_ _0047_ clknet_4_9_0_Clock B\[1\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5814_ _3026_ _0980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6794_ _1914_ _1921_ _1922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_37_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8533_ _0088_ _3681_ _3728_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5745_ _0867_ _0887_ _0917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8464_ net14 _3663_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5676_ _0802_ _0847_ _0848_ _0849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8161__A1 _3261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7415_ _2511_ _2512_ _2559_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4627_ B\[1\]\[5\] _3780_ _3271_ _3783_ _3949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_117_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8395_ _3592_ _3595_ _3596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_1350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6711__A2 _1841_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4558_ _3852_ _3879_ _3881_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_11_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7346_ _3874_ _1952_ _2485_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4489_ A\[2\]\[0\] _3744_ _3391_ _3750_ _3701_ _3812_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_7277_ _0980_ _2101_ _2410_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6228_ _4161_ _0038_ _1381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8216__A2 _2152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6159_ _1164_ _0044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5450__A2 _0390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7727__A1 C\[0\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6950__A2 _2001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4713__A1 B\[3\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4713__B2 _2919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7663__B1 _1972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6218__A1 _1372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7718__A1 _0348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7718__B2 _2872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5530_ _0701_ _0706_ _0707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4952__A1 _4263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4689__I _3830_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5461_ _3805_ _0487_ _0638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4412_ _3174_ _3337_ _3662_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7200_ _2252_ _2263_ _2326_ _2327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5392_ _0568_ _0569_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8180_ _3286_ _3364_ _3365_ _3366_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7131_ _2138_ _2249_ _2251_ _2252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4343_ _2298_ _2930_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7062_ _3960_ _3861_ _1755_ _2183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_99_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6013_ _3993_ _3790_ _4093_ _1027_ _1176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_101_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7957__A1 _0822_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7964_ _3099_ _3134_ _3135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_55_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5432__A2 _0529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6915_ _2029_ _2037_ _2038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_74_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4373__B A\[3\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7895_ _2979_ _2988_ _3059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7709__A1 _0761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6846_ _1971_ _1972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8509__I0 _0097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6777_ _1905_ _1906_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8516_ _0129_ _3670_ _3712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5728_ _0774_ _0899_ _0900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8134__A1 _0647_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4599__I _3920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8447_ C\[0\]\[15\] _3462_ _0007_ _3600_ _3651_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_5659_ _0827_ _0830_ _0832_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6696__A1 _1824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8378_ _3508_ _3532_ _3578_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_105_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7329_ _2385_ _2451_ _2465_ _2466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6448__A1 _0031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5671__A2 _0498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7948__A1 _3018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8681__D _0074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5423__A2 _0582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6620__A1 _1753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5187__A1 _4071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6923__A2 _2045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8125__A1 _3305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer6 _1889_ net39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
XANTENNA__4302__I _2383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5111__A1 _0285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5133__I _0314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5662__A2 _0834_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4465__A3 _2513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8591__D _0036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4961_ _3965_ _4275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6700_ _3962_ _1772_ _1832_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7680_ _2792_ _2833_ _2834_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4892_ _4207_ _0028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8364__A1 _3553_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5178__A1 _3456_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6631_ _4116_ _1703_ _1749_ _1765_ _1766_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__4925__A1 C\[3\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6562_ _1701_ _1702_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8301_ _3378_ _3496_ _3447_ _3448_ _3497_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5513_ _0686_ _0688_ _0690_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6493_ _1635_ _1636_ _1637_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8232_ _3344_ _3346_ _3419_ _3422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5444_ _0606_ _0620_ _0621_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_12_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8163_ _3344_ _3346_ _3348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5375_ _0549_ _0550_ _0551_ _0552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7114_ _3861_ _1808_ _2235_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4326_ _2394_ _2755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_113_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8094_ _3198_ _3235_ _3273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7045_ _2160_ _2162_ _2165_ _2166_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_80_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5653__A2 _3871_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4882__I _3848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8052__B1 _1732_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7947_ _3019_ _1980_ _3116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7878_ _2970_ _3042_ _3043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8355__A1 _3518_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6829_ _1945_ _1954_ _1955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_23_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6602__I _1700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8107__A1 _0577_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5184__A4 _0355_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7330__A2 _2391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8676__D _0083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7433__I _2123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6841__A1 _4200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4792__I _2438_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7608__I _0467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5580__A1 _3822_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5128__I _4031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8586__D _0031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7872__A3 _3035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5160_ _0309_ _0322_ _0341_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_116_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5091_ _0267_ _0269_ _0273_ _0274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_110_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7624__A3 _2776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7388__A2 _2462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7801_ _2921_ _2924_ _2960_ _2961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_77_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5399__A1 _3894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5399__B2 B\[2\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5993_ _1152_ _1155_ _1156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_91_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7732_ _2858_ _2887_ _2888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4944_ _4256_ _4257_ _4259_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_80_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4610__A3 _3921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7663_ _2815_ _1771_ _1972_ _2773_ _2817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4875_ _4120_ _4191_ _4192_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_127_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6614_ _1738_ _1750_ _1751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7594_ _2744_ _2746_ _2747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_118_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6545_ _1656_ _1660_ _1684_ _1685_ _1686_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4374__A2 net10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6476_ _1400_ _1404_ _1620_ _1554_ _1621_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_106_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8215_ _3397_ _3404_ _3405_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5427_ _0532_ _0602_ _0603_ _0604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5874__A2 _1038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8146_ _3270_ _3329_ _3330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5358_ _3806_ _0398_ _0413_ _0533_ _0535_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_114_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4309_ _2567_ _2578_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_102_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8077_ _3160_ _3166_ _3254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5289_ _0466_ _0467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7028_ _1985_ _1907_ _2149_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4834__B1 _3894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4601__A3 _3817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7000__A1 _4113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7551__A2 _0947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4365__A2 _3144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5562__A1 _0512_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8500__A1 _3696_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7303__A2 _2437_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4787__I _3899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5314__A1 _0489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5865__A2 _4067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7067__A1 _2178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6290__A2 _3981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8319__A1 _0481_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7790__A2 _3929_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8573__CLK clknet_4_3_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4660_ _3890_ _3982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5553__A1 _0629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4591_ _3885_ _3886_ _3913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_143_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6330_ _1479_ C\[2\]\[13\] _0469_ _1480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6261_ _1305_ _1331_ _1412_ _1413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8000_ _3169_ _3170_ _3171_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5212_ _0392_ _0393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6192_ _1228_ _1237_ _1348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5143_ net44 _0304_ _0306_ B\[2\]\[6\] _0325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_96_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5608__A2 _0370_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5074_ _0234_ _0252_ _0257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5321__I _0461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7230__A1 _1985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5976_ _1012_ _0989_ _1042_ _1139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7781__A2 _0352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7715_ _2868_ _2822_ _2869_ _2870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4927_ _3927_ _4242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8695_ _0141_ clknet_4_7_0_Clock net31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7646_ _2761_ _0011_ _2797_ _2798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4858_ _4171_ _4174_ _4175_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_53_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4347__A2 _2963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5544__A1 _4169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7577_ _2731_ _0094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4789_ _4106_ _4108_ _4109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_88_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6528_ _1583_ _1643_ _1668_ _1588_ _1669_ _1670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_118_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7297__A1 _2364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6459_ _1527_ _1540_ _1604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_109_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5847__A2 _4188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4400__I _3531_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8129_ _3309_ _3231_ _3310_ _3311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_76_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4283__A1 _2233_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8549__A1 _3737_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7867__B _3030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8013__A3 _2050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8596__CLK clknet_4_3_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7772__A2 _2928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5387__B B\[0\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7158__I _2281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5535__A1 _3973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8485__B1 _3684_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5299__B1 _0474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5838__A2 _1002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4510__A2 _3832_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6263__A2 _3900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7460__A1 _2602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5830_ _0994_ _0995_ _0996_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7763__A2 _2918_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5761_ _0928_ _0929_ _0931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7500_ _2636_ _2649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4712_ _3858_ _4033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8480_ _3678_ _0094_ _3679_ _3680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5692_ _0817_ _0818_ _0865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7431_ _2510_ _2574_ _2575_ _2514_ _2509_ _2576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_4643_ _3964_ _3965_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7362_ _4069_ _1529_ _0004_ _2501_ _2502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4574_ _3891_ _3895_ _3821_ _3896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7279__A1 _0060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6313_ _1349_ _1353_ _1463_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7279__B2 _0059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7293_ _2423_ _2426_ _2428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5316__I _0376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6244_ _1394_ _1396_ _1397_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6856__B A\[0\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6175_ _1305_ _1331_ _1332_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_58_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5126_ _0307_ _0308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5057_ _0193_ _0194_ _0240_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_72_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7203__A1 _2313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6006__A2 _1029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7754__A2 _2865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5765__A1 _0919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5959_ _1122_ _1123_ _1124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8678_ _0085_ clknet_4_7_0_Clock C\[3\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5517__A1 _0625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7629_ _2766_ _2781_ _2782_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_103_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6610__I _1746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4740__A2 _3769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8537__I _3730_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8684__D _0077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7442__A1 _2536_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5756__A1 _0024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8170__A2 _3294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8611__CLK clknet_4_1_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5136__I _0317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4290_ _2362_ _2373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_125_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5287__A3 _0464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8594__D _0039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7980_ _3149_ _0129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7984__A2 _3135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6931_ _1998_ _2054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_78_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6862_ _1986_ _1987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8601_ _0046_ clknet_4_3_0_Clock B\[1\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5813_ _4124_ _4145_ _0979_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6793_ _1915_ _1920_ _1921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8532_ _3692_ _3725_ _3708_ _3726_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5744_ _0914_ _0915_ _0916_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_124_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8536__I1 _0074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8463_ _3661_ _3796_ _0019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5675_ _0799_ _0844_ _0848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7414_ _2550_ _2551_ _2557_ _2558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_129_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4626_ _3947_ _3948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8394_ _3500_ _3594_ _3595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6711__A3 _1842_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7345_ _3877_ _2123_ _2484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4557_ _3852_ _3879_ _3880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5046__I _0222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7276_ _2403_ _2408_ _2409_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4488_ _3758_ _3774_ _3801_ _3810_ _3811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_132_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7672__A1 _0035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6227_ _0718_ _0038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6158_ _0045_ _4161_ _1316_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5109_ _0281_ _0290_ _0292_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_57_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6089_ _0419_ _0658_ _1248_ _0468_ _1250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_3427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5435__B1 _0355_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7188__B1 _2229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7727__A2 _4239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8634__CLK clknet_4_11_0_Clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8679__D _0086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6163__A1 _3794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4713__A2 _2930_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5910__A1 _0704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput30 net30 Result[7] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_107_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4795__I _3326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7663__A1 _2815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7663__B2 _2773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4477__A1 _3794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6218__A2 C\[2\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7718__A2 _0352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8391__A2 _0015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4401__A1 _3542_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8589__D _0034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4952__A2 _4264_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8143__A2 _3325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5460_ _0574_ _0493_ _0637_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4411_ _3646_ _0030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5391_ _0504_ _0505_ _3593_ _0568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7130_ _0043_ _2250_ _2141_ _2251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4342_ _2908_ _2919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_82_1508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7061_ _2051_ _2180_ _2181_ _2182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__8177__I _3289_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4468__A1 _3778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6012_ _1172_ _1173_ _1174_ _1175_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_113_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
.ends

