magic
tech gf180mcuC
magscale 1 5
timestamp 1670203860
<< obsm1 >>
rect 672 855 199304 148273
<< metal2 >>
rect 1848 149600 1904 150000
rect 3584 149600 3640 150000
rect 5320 149600 5376 150000
rect 7056 149600 7112 150000
rect 8792 149600 8848 150000
rect 10528 149600 10584 150000
rect 12264 149600 12320 150000
rect 14000 149600 14056 150000
rect 15736 149600 15792 150000
rect 17472 149600 17528 150000
rect 19208 149600 19264 150000
rect 20944 149600 21000 150000
rect 22680 149600 22736 150000
rect 24416 149600 24472 150000
rect 26152 149600 26208 150000
rect 27888 149600 27944 150000
rect 29624 149600 29680 150000
rect 31360 149600 31416 150000
rect 33096 149600 33152 150000
rect 34832 149600 34888 150000
rect 36568 149600 36624 150000
rect 38304 149600 38360 150000
rect 40040 149600 40096 150000
rect 41776 149600 41832 150000
rect 43512 149600 43568 150000
rect 45248 149600 45304 150000
rect 46984 149600 47040 150000
rect 48720 149600 48776 150000
rect 50456 149600 50512 150000
rect 52192 149600 52248 150000
rect 53928 149600 53984 150000
rect 55664 149600 55720 150000
rect 57400 149600 57456 150000
rect 59136 149600 59192 150000
rect 60872 149600 60928 150000
rect 62608 149600 62664 150000
rect 64344 149600 64400 150000
rect 66080 149600 66136 150000
rect 67816 149600 67872 150000
rect 69552 149600 69608 150000
rect 71288 149600 71344 150000
rect 73024 149600 73080 150000
rect 74760 149600 74816 150000
rect 76496 149600 76552 150000
rect 78232 149600 78288 150000
rect 79968 149600 80024 150000
rect 81704 149600 81760 150000
rect 83440 149600 83496 150000
rect 85176 149600 85232 150000
rect 86912 149600 86968 150000
rect 88648 149600 88704 150000
rect 90384 149600 90440 150000
rect 92120 149600 92176 150000
rect 93856 149600 93912 150000
rect 95592 149600 95648 150000
rect 97328 149600 97384 150000
rect 99064 149600 99120 150000
rect 100800 149600 100856 150000
rect 102536 149600 102592 150000
rect 104272 149600 104328 150000
rect 106008 149600 106064 150000
rect 107744 149600 107800 150000
rect 109480 149600 109536 150000
rect 111216 149600 111272 150000
rect 112952 149600 113008 150000
rect 114688 149600 114744 150000
rect 116424 149600 116480 150000
rect 118160 149600 118216 150000
rect 119896 149600 119952 150000
rect 121632 149600 121688 150000
rect 123368 149600 123424 150000
rect 125104 149600 125160 150000
rect 126840 149600 126896 150000
rect 128576 149600 128632 150000
rect 130312 149600 130368 150000
rect 132048 149600 132104 150000
rect 133784 149600 133840 150000
rect 135520 149600 135576 150000
rect 137256 149600 137312 150000
rect 138992 149600 139048 150000
rect 140728 149600 140784 150000
rect 142464 149600 142520 150000
rect 144200 149600 144256 150000
rect 145936 149600 145992 150000
rect 147672 149600 147728 150000
rect 149408 149600 149464 150000
rect 151144 149600 151200 150000
rect 152880 149600 152936 150000
rect 154616 149600 154672 150000
rect 156352 149600 156408 150000
rect 158088 149600 158144 150000
rect 159824 149600 159880 150000
rect 161560 149600 161616 150000
rect 163296 149600 163352 150000
rect 165032 149600 165088 150000
rect 166768 149600 166824 150000
rect 168504 149600 168560 150000
rect 170240 149600 170296 150000
rect 171976 149600 172032 150000
rect 173712 149600 173768 150000
rect 175448 149600 175504 150000
rect 177184 149600 177240 150000
rect 178920 149600 178976 150000
rect 180656 149600 180712 150000
rect 182392 149600 182448 150000
rect 184128 149600 184184 150000
rect 185864 149600 185920 150000
rect 187600 149600 187656 150000
rect 189336 149600 189392 150000
rect 191072 149600 191128 150000
rect 192808 149600 192864 150000
rect 194544 149600 194600 150000
rect 196280 149600 196336 150000
rect 198016 149600 198072 150000
rect 3528 0 3584 400
rect 3920 0 3976 400
rect 4312 0 4368 400
rect 4704 0 4760 400
rect 5096 0 5152 400
rect 5488 0 5544 400
rect 5880 0 5936 400
rect 6272 0 6328 400
rect 6664 0 6720 400
rect 7056 0 7112 400
rect 7448 0 7504 400
rect 7840 0 7896 400
rect 8232 0 8288 400
rect 8624 0 8680 400
rect 9016 0 9072 400
rect 9408 0 9464 400
rect 9800 0 9856 400
rect 10192 0 10248 400
rect 10584 0 10640 400
rect 10976 0 11032 400
rect 11368 0 11424 400
rect 11760 0 11816 400
rect 12152 0 12208 400
rect 12544 0 12600 400
rect 12936 0 12992 400
rect 13328 0 13384 400
rect 13720 0 13776 400
rect 14112 0 14168 400
rect 14504 0 14560 400
rect 14896 0 14952 400
rect 15288 0 15344 400
rect 15680 0 15736 400
rect 16072 0 16128 400
rect 16464 0 16520 400
rect 16856 0 16912 400
rect 17248 0 17304 400
rect 17640 0 17696 400
rect 18032 0 18088 400
rect 18424 0 18480 400
rect 18816 0 18872 400
rect 19208 0 19264 400
rect 19600 0 19656 400
rect 19992 0 20048 400
rect 20384 0 20440 400
rect 20776 0 20832 400
rect 21168 0 21224 400
rect 21560 0 21616 400
rect 21952 0 22008 400
rect 22344 0 22400 400
rect 22736 0 22792 400
rect 23128 0 23184 400
rect 23520 0 23576 400
rect 23912 0 23968 400
rect 24304 0 24360 400
rect 24696 0 24752 400
rect 25088 0 25144 400
rect 25480 0 25536 400
rect 25872 0 25928 400
rect 26264 0 26320 400
rect 26656 0 26712 400
rect 27048 0 27104 400
rect 27440 0 27496 400
rect 27832 0 27888 400
rect 28224 0 28280 400
rect 28616 0 28672 400
rect 29008 0 29064 400
rect 29400 0 29456 400
rect 29792 0 29848 400
rect 30184 0 30240 400
rect 30576 0 30632 400
rect 30968 0 31024 400
rect 31360 0 31416 400
rect 31752 0 31808 400
rect 32144 0 32200 400
rect 32536 0 32592 400
rect 32928 0 32984 400
rect 33320 0 33376 400
rect 33712 0 33768 400
rect 34104 0 34160 400
rect 34496 0 34552 400
rect 34888 0 34944 400
rect 35280 0 35336 400
rect 35672 0 35728 400
rect 36064 0 36120 400
rect 36456 0 36512 400
rect 36848 0 36904 400
rect 37240 0 37296 400
rect 37632 0 37688 400
rect 38024 0 38080 400
rect 38416 0 38472 400
rect 38808 0 38864 400
rect 39200 0 39256 400
rect 39592 0 39648 400
rect 39984 0 40040 400
rect 40376 0 40432 400
rect 40768 0 40824 400
rect 41160 0 41216 400
rect 41552 0 41608 400
rect 41944 0 42000 400
rect 42336 0 42392 400
rect 42728 0 42784 400
rect 43120 0 43176 400
rect 43512 0 43568 400
rect 43904 0 43960 400
rect 44296 0 44352 400
rect 44688 0 44744 400
rect 45080 0 45136 400
rect 45472 0 45528 400
rect 45864 0 45920 400
rect 46256 0 46312 400
rect 46648 0 46704 400
rect 47040 0 47096 400
rect 47432 0 47488 400
rect 47824 0 47880 400
rect 48216 0 48272 400
rect 48608 0 48664 400
rect 49000 0 49056 400
rect 49392 0 49448 400
rect 49784 0 49840 400
rect 50176 0 50232 400
rect 50568 0 50624 400
rect 50960 0 51016 400
rect 51352 0 51408 400
rect 51744 0 51800 400
rect 52136 0 52192 400
rect 52528 0 52584 400
rect 52920 0 52976 400
rect 53312 0 53368 400
rect 53704 0 53760 400
rect 54096 0 54152 400
rect 54488 0 54544 400
rect 54880 0 54936 400
rect 55272 0 55328 400
rect 55664 0 55720 400
rect 56056 0 56112 400
rect 56448 0 56504 400
rect 56840 0 56896 400
rect 57232 0 57288 400
rect 57624 0 57680 400
rect 58016 0 58072 400
rect 58408 0 58464 400
rect 58800 0 58856 400
rect 59192 0 59248 400
rect 59584 0 59640 400
rect 59976 0 60032 400
rect 60368 0 60424 400
rect 60760 0 60816 400
rect 61152 0 61208 400
rect 61544 0 61600 400
rect 61936 0 61992 400
rect 62328 0 62384 400
rect 62720 0 62776 400
rect 63112 0 63168 400
rect 63504 0 63560 400
rect 63896 0 63952 400
rect 64288 0 64344 400
rect 64680 0 64736 400
rect 65072 0 65128 400
rect 65464 0 65520 400
rect 65856 0 65912 400
rect 66248 0 66304 400
rect 66640 0 66696 400
rect 67032 0 67088 400
rect 67424 0 67480 400
rect 67816 0 67872 400
rect 68208 0 68264 400
rect 68600 0 68656 400
rect 68992 0 69048 400
rect 69384 0 69440 400
rect 69776 0 69832 400
rect 70168 0 70224 400
rect 70560 0 70616 400
rect 70952 0 71008 400
rect 71344 0 71400 400
rect 71736 0 71792 400
rect 72128 0 72184 400
rect 72520 0 72576 400
rect 72912 0 72968 400
rect 73304 0 73360 400
rect 73696 0 73752 400
rect 74088 0 74144 400
rect 74480 0 74536 400
rect 74872 0 74928 400
rect 75264 0 75320 400
rect 75656 0 75712 400
rect 76048 0 76104 400
rect 76440 0 76496 400
rect 76832 0 76888 400
rect 77224 0 77280 400
rect 77616 0 77672 400
rect 78008 0 78064 400
rect 78400 0 78456 400
rect 78792 0 78848 400
rect 79184 0 79240 400
rect 79576 0 79632 400
rect 79968 0 80024 400
rect 80360 0 80416 400
rect 80752 0 80808 400
rect 81144 0 81200 400
rect 81536 0 81592 400
rect 81928 0 81984 400
rect 82320 0 82376 400
rect 82712 0 82768 400
rect 83104 0 83160 400
rect 83496 0 83552 400
rect 83888 0 83944 400
rect 84280 0 84336 400
rect 84672 0 84728 400
rect 85064 0 85120 400
rect 85456 0 85512 400
rect 85848 0 85904 400
rect 86240 0 86296 400
rect 86632 0 86688 400
rect 87024 0 87080 400
rect 87416 0 87472 400
rect 87808 0 87864 400
rect 88200 0 88256 400
rect 88592 0 88648 400
rect 88984 0 89040 400
rect 89376 0 89432 400
rect 89768 0 89824 400
rect 90160 0 90216 400
rect 90552 0 90608 400
rect 90944 0 91000 400
rect 91336 0 91392 400
rect 91728 0 91784 400
rect 92120 0 92176 400
rect 92512 0 92568 400
rect 92904 0 92960 400
rect 93296 0 93352 400
rect 93688 0 93744 400
rect 94080 0 94136 400
rect 94472 0 94528 400
rect 94864 0 94920 400
rect 95256 0 95312 400
rect 95648 0 95704 400
rect 96040 0 96096 400
rect 96432 0 96488 400
rect 96824 0 96880 400
rect 97216 0 97272 400
rect 97608 0 97664 400
rect 98000 0 98056 400
rect 98392 0 98448 400
rect 98784 0 98840 400
rect 99176 0 99232 400
rect 99568 0 99624 400
rect 99960 0 100016 400
rect 100352 0 100408 400
rect 100744 0 100800 400
rect 101136 0 101192 400
rect 101528 0 101584 400
rect 101920 0 101976 400
rect 102312 0 102368 400
rect 102704 0 102760 400
rect 103096 0 103152 400
rect 103488 0 103544 400
rect 103880 0 103936 400
rect 104272 0 104328 400
rect 104664 0 104720 400
rect 105056 0 105112 400
rect 105448 0 105504 400
rect 105840 0 105896 400
rect 106232 0 106288 400
rect 106624 0 106680 400
rect 107016 0 107072 400
rect 107408 0 107464 400
rect 107800 0 107856 400
rect 108192 0 108248 400
rect 108584 0 108640 400
rect 108976 0 109032 400
rect 109368 0 109424 400
rect 109760 0 109816 400
rect 110152 0 110208 400
rect 110544 0 110600 400
rect 110936 0 110992 400
rect 111328 0 111384 400
rect 111720 0 111776 400
rect 112112 0 112168 400
rect 112504 0 112560 400
rect 112896 0 112952 400
rect 113288 0 113344 400
rect 113680 0 113736 400
rect 114072 0 114128 400
rect 114464 0 114520 400
rect 114856 0 114912 400
rect 115248 0 115304 400
rect 115640 0 115696 400
rect 116032 0 116088 400
rect 116424 0 116480 400
rect 116816 0 116872 400
rect 117208 0 117264 400
rect 117600 0 117656 400
rect 117992 0 118048 400
rect 118384 0 118440 400
rect 118776 0 118832 400
rect 119168 0 119224 400
rect 119560 0 119616 400
rect 119952 0 120008 400
rect 120344 0 120400 400
rect 120736 0 120792 400
rect 121128 0 121184 400
rect 121520 0 121576 400
rect 121912 0 121968 400
rect 122304 0 122360 400
rect 122696 0 122752 400
rect 123088 0 123144 400
rect 123480 0 123536 400
rect 123872 0 123928 400
rect 124264 0 124320 400
rect 124656 0 124712 400
rect 125048 0 125104 400
rect 125440 0 125496 400
rect 125832 0 125888 400
rect 126224 0 126280 400
rect 126616 0 126672 400
rect 127008 0 127064 400
rect 127400 0 127456 400
rect 127792 0 127848 400
rect 128184 0 128240 400
rect 128576 0 128632 400
rect 128968 0 129024 400
rect 129360 0 129416 400
rect 129752 0 129808 400
rect 130144 0 130200 400
rect 130536 0 130592 400
rect 130928 0 130984 400
rect 131320 0 131376 400
rect 131712 0 131768 400
rect 132104 0 132160 400
rect 132496 0 132552 400
rect 132888 0 132944 400
rect 133280 0 133336 400
rect 133672 0 133728 400
rect 134064 0 134120 400
rect 134456 0 134512 400
rect 134848 0 134904 400
rect 135240 0 135296 400
rect 135632 0 135688 400
rect 136024 0 136080 400
rect 136416 0 136472 400
rect 136808 0 136864 400
rect 137200 0 137256 400
rect 137592 0 137648 400
rect 137984 0 138040 400
rect 138376 0 138432 400
rect 138768 0 138824 400
rect 139160 0 139216 400
rect 139552 0 139608 400
rect 139944 0 140000 400
rect 140336 0 140392 400
rect 140728 0 140784 400
rect 141120 0 141176 400
rect 141512 0 141568 400
rect 141904 0 141960 400
rect 142296 0 142352 400
rect 142688 0 142744 400
rect 143080 0 143136 400
rect 143472 0 143528 400
rect 143864 0 143920 400
rect 144256 0 144312 400
rect 144648 0 144704 400
rect 145040 0 145096 400
rect 145432 0 145488 400
rect 145824 0 145880 400
rect 146216 0 146272 400
rect 146608 0 146664 400
rect 147000 0 147056 400
rect 147392 0 147448 400
rect 147784 0 147840 400
rect 148176 0 148232 400
rect 148568 0 148624 400
rect 148960 0 149016 400
rect 149352 0 149408 400
rect 149744 0 149800 400
rect 150136 0 150192 400
rect 150528 0 150584 400
rect 150920 0 150976 400
rect 151312 0 151368 400
rect 151704 0 151760 400
rect 152096 0 152152 400
rect 152488 0 152544 400
rect 152880 0 152936 400
rect 153272 0 153328 400
rect 153664 0 153720 400
rect 154056 0 154112 400
rect 154448 0 154504 400
rect 154840 0 154896 400
rect 155232 0 155288 400
rect 155624 0 155680 400
rect 156016 0 156072 400
rect 156408 0 156464 400
rect 156800 0 156856 400
rect 157192 0 157248 400
rect 157584 0 157640 400
rect 157976 0 158032 400
rect 158368 0 158424 400
rect 158760 0 158816 400
rect 159152 0 159208 400
rect 159544 0 159600 400
rect 159936 0 159992 400
rect 160328 0 160384 400
rect 160720 0 160776 400
rect 161112 0 161168 400
rect 161504 0 161560 400
rect 161896 0 161952 400
rect 162288 0 162344 400
rect 162680 0 162736 400
rect 163072 0 163128 400
rect 163464 0 163520 400
rect 163856 0 163912 400
rect 164248 0 164304 400
rect 164640 0 164696 400
rect 165032 0 165088 400
rect 165424 0 165480 400
rect 165816 0 165872 400
rect 166208 0 166264 400
rect 166600 0 166656 400
rect 166992 0 167048 400
rect 167384 0 167440 400
rect 167776 0 167832 400
rect 168168 0 168224 400
rect 168560 0 168616 400
rect 168952 0 169008 400
rect 169344 0 169400 400
rect 169736 0 169792 400
rect 170128 0 170184 400
rect 170520 0 170576 400
rect 170912 0 170968 400
rect 171304 0 171360 400
rect 171696 0 171752 400
rect 172088 0 172144 400
rect 172480 0 172536 400
rect 172872 0 172928 400
rect 173264 0 173320 400
rect 173656 0 173712 400
rect 174048 0 174104 400
rect 174440 0 174496 400
rect 174832 0 174888 400
rect 175224 0 175280 400
rect 175616 0 175672 400
rect 176008 0 176064 400
rect 176400 0 176456 400
rect 176792 0 176848 400
rect 177184 0 177240 400
rect 177576 0 177632 400
rect 177968 0 178024 400
rect 178360 0 178416 400
rect 178752 0 178808 400
rect 179144 0 179200 400
rect 179536 0 179592 400
rect 179928 0 179984 400
rect 180320 0 180376 400
rect 180712 0 180768 400
rect 181104 0 181160 400
rect 181496 0 181552 400
rect 181888 0 181944 400
rect 182280 0 182336 400
rect 182672 0 182728 400
rect 183064 0 183120 400
rect 183456 0 183512 400
rect 183848 0 183904 400
rect 184240 0 184296 400
rect 184632 0 184688 400
rect 185024 0 185080 400
rect 185416 0 185472 400
rect 185808 0 185864 400
rect 186200 0 186256 400
rect 186592 0 186648 400
rect 186984 0 187040 400
rect 187376 0 187432 400
rect 187768 0 187824 400
rect 188160 0 188216 400
rect 188552 0 188608 400
rect 188944 0 189000 400
rect 189336 0 189392 400
rect 189728 0 189784 400
rect 190120 0 190176 400
rect 190512 0 190568 400
rect 190904 0 190960 400
rect 191296 0 191352 400
rect 191688 0 191744 400
rect 192080 0 192136 400
rect 192472 0 192528 400
rect 192864 0 192920 400
rect 193256 0 193312 400
rect 193648 0 193704 400
rect 194040 0 194096 400
rect 194432 0 194488 400
rect 194824 0 194880 400
rect 195216 0 195272 400
rect 195608 0 195664 400
rect 196000 0 196056 400
rect 196392 0 196448 400
<< obsm2 >>
rect 2238 149570 3554 149600
rect 3670 149570 5290 149600
rect 5406 149570 7026 149600
rect 7142 149570 8762 149600
rect 8878 149570 10498 149600
rect 10614 149570 12234 149600
rect 12350 149570 13970 149600
rect 14086 149570 15706 149600
rect 15822 149570 17442 149600
rect 17558 149570 19178 149600
rect 19294 149570 20914 149600
rect 21030 149570 22650 149600
rect 22766 149570 24386 149600
rect 24502 149570 26122 149600
rect 26238 149570 27858 149600
rect 27974 149570 29594 149600
rect 29710 149570 31330 149600
rect 31446 149570 33066 149600
rect 33182 149570 34802 149600
rect 34918 149570 36538 149600
rect 36654 149570 38274 149600
rect 38390 149570 40010 149600
rect 40126 149570 41746 149600
rect 41862 149570 43482 149600
rect 43598 149570 45218 149600
rect 45334 149570 46954 149600
rect 47070 149570 48690 149600
rect 48806 149570 50426 149600
rect 50542 149570 52162 149600
rect 52278 149570 53898 149600
rect 54014 149570 55634 149600
rect 55750 149570 57370 149600
rect 57486 149570 59106 149600
rect 59222 149570 60842 149600
rect 60958 149570 62578 149600
rect 62694 149570 64314 149600
rect 64430 149570 66050 149600
rect 66166 149570 67786 149600
rect 67902 149570 69522 149600
rect 69638 149570 71258 149600
rect 71374 149570 72994 149600
rect 73110 149570 74730 149600
rect 74846 149570 76466 149600
rect 76582 149570 78202 149600
rect 78318 149570 79938 149600
rect 80054 149570 81674 149600
rect 81790 149570 83410 149600
rect 83526 149570 85146 149600
rect 85262 149570 86882 149600
rect 86998 149570 88618 149600
rect 88734 149570 90354 149600
rect 90470 149570 92090 149600
rect 92206 149570 93826 149600
rect 93942 149570 95562 149600
rect 95678 149570 97298 149600
rect 97414 149570 99034 149600
rect 99150 149570 100770 149600
rect 100886 149570 102506 149600
rect 102622 149570 104242 149600
rect 104358 149570 105978 149600
rect 106094 149570 107714 149600
rect 107830 149570 109450 149600
rect 109566 149570 111186 149600
rect 111302 149570 112922 149600
rect 113038 149570 114658 149600
rect 114774 149570 116394 149600
rect 116510 149570 118130 149600
rect 118246 149570 119866 149600
rect 119982 149570 121602 149600
rect 121718 149570 123338 149600
rect 123454 149570 125074 149600
rect 125190 149570 126810 149600
rect 126926 149570 128546 149600
rect 128662 149570 130282 149600
rect 130398 149570 132018 149600
rect 132134 149570 133754 149600
rect 133870 149570 135490 149600
rect 135606 149570 137226 149600
rect 137342 149570 138962 149600
rect 139078 149570 140698 149600
rect 140814 149570 142434 149600
rect 142550 149570 144170 149600
rect 144286 149570 145906 149600
rect 146022 149570 147642 149600
rect 147758 149570 149378 149600
rect 149494 149570 151114 149600
rect 151230 149570 152850 149600
rect 152966 149570 154586 149600
rect 154702 149570 156322 149600
rect 156438 149570 158058 149600
rect 158174 149570 159794 149600
rect 159910 149570 161530 149600
rect 161646 149570 163266 149600
rect 163382 149570 165002 149600
rect 165118 149570 166738 149600
rect 166854 149570 168474 149600
rect 168590 149570 170210 149600
rect 170326 149570 171946 149600
rect 172062 149570 173682 149600
rect 173798 149570 175418 149600
rect 175534 149570 177154 149600
rect 177270 149570 178890 149600
rect 179006 149570 180626 149600
rect 180742 149570 182362 149600
rect 182478 149570 184098 149600
rect 184214 149570 185834 149600
rect 185950 149570 187570 149600
rect 187686 149570 189306 149600
rect 189422 149570 191042 149600
rect 191158 149570 192778 149600
rect 192894 149570 194514 149600
rect 194630 149570 196250 149600
rect 196366 149570 197986 149600
rect 198102 149570 198170 149600
rect 2238 430 198170 149570
rect 2238 400 3498 430
rect 3614 400 3890 430
rect 4006 400 4282 430
rect 4398 400 4674 430
rect 4790 400 5066 430
rect 5182 400 5458 430
rect 5574 400 5850 430
rect 5966 400 6242 430
rect 6358 400 6634 430
rect 6750 400 7026 430
rect 7142 400 7418 430
rect 7534 400 7810 430
rect 7926 400 8202 430
rect 8318 400 8594 430
rect 8710 400 8986 430
rect 9102 400 9378 430
rect 9494 400 9770 430
rect 9886 400 10162 430
rect 10278 400 10554 430
rect 10670 400 10946 430
rect 11062 400 11338 430
rect 11454 400 11730 430
rect 11846 400 12122 430
rect 12238 400 12514 430
rect 12630 400 12906 430
rect 13022 400 13298 430
rect 13414 400 13690 430
rect 13806 400 14082 430
rect 14198 400 14474 430
rect 14590 400 14866 430
rect 14982 400 15258 430
rect 15374 400 15650 430
rect 15766 400 16042 430
rect 16158 400 16434 430
rect 16550 400 16826 430
rect 16942 400 17218 430
rect 17334 400 17610 430
rect 17726 400 18002 430
rect 18118 400 18394 430
rect 18510 400 18786 430
rect 18902 400 19178 430
rect 19294 400 19570 430
rect 19686 400 19962 430
rect 20078 400 20354 430
rect 20470 400 20746 430
rect 20862 400 21138 430
rect 21254 400 21530 430
rect 21646 400 21922 430
rect 22038 400 22314 430
rect 22430 400 22706 430
rect 22822 400 23098 430
rect 23214 400 23490 430
rect 23606 400 23882 430
rect 23998 400 24274 430
rect 24390 400 24666 430
rect 24782 400 25058 430
rect 25174 400 25450 430
rect 25566 400 25842 430
rect 25958 400 26234 430
rect 26350 400 26626 430
rect 26742 400 27018 430
rect 27134 400 27410 430
rect 27526 400 27802 430
rect 27918 400 28194 430
rect 28310 400 28586 430
rect 28702 400 28978 430
rect 29094 400 29370 430
rect 29486 400 29762 430
rect 29878 400 30154 430
rect 30270 400 30546 430
rect 30662 400 30938 430
rect 31054 400 31330 430
rect 31446 400 31722 430
rect 31838 400 32114 430
rect 32230 400 32506 430
rect 32622 400 32898 430
rect 33014 400 33290 430
rect 33406 400 33682 430
rect 33798 400 34074 430
rect 34190 400 34466 430
rect 34582 400 34858 430
rect 34974 400 35250 430
rect 35366 400 35642 430
rect 35758 400 36034 430
rect 36150 400 36426 430
rect 36542 400 36818 430
rect 36934 400 37210 430
rect 37326 400 37602 430
rect 37718 400 37994 430
rect 38110 400 38386 430
rect 38502 400 38778 430
rect 38894 400 39170 430
rect 39286 400 39562 430
rect 39678 400 39954 430
rect 40070 400 40346 430
rect 40462 400 40738 430
rect 40854 400 41130 430
rect 41246 400 41522 430
rect 41638 400 41914 430
rect 42030 400 42306 430
rect 42422 400 42698 430
rect 42814 400 43090 430
rect 43206 400 43482 430
rect 43598 400 43874 430
rect 43990 400 44266 430
rect 44382 400 44658 430
rect 44774 400 45050 430
rect 45166 400 45442 430
rect 45558 400 45834 430
rect 45950 400 46226 430
rect 46342 400 46618 430
rect 46734 400 47010 430
rect 47126 400 47402 430
rect 47518 400 47794 430
rect 47910 400 48186 430
rect 48302 400 48578 430
rect 48694 400 48970 430
rect 49086 400 49362 430
rect 49478 400 49754 430
rect 49870 400 50146 430
rect 50262 400 50538 430
rect 50654 400 50930 430
rect 51046 400 51322 430
rect 51438 400 51714 430
rect 51830 400 52106 430
rect 52222 400 52498 430
rect 52614 400 52890 430
rect 53006 400 53282 430
rect 53398 400 53674 430
rect 53790 400 54066 430
rect 54182 400 54458 430
rect 54574 400 54850 430
rect 54966 400 55242 430
rect 55358 400 55634 430
rect 55750 400 56026 430
rect 56142 400 56418 430
rect 56534 400 56810 430
rect 56926 400 57202 430
rect 57318 400 57594 430
rect 57710 400 57986 430
rect 58102 400 58378 430
rect 58494 400 58770 430
rect 58886 400 59162 430
rect 59278 400 59554 430
rect 59670 400 59946 430
rect 60062 400 60338 430
rect 60454 400 60730 430
rect 60846 400 61122 430
rect 61238 400 61514 430
rect 61630 400 61906 430
rect 62022 400 62298 430
rect 62414 400 62690 430
rect 62806 400 63082 430
rect 63198 400 63474 430
rect 63590 400 63866 430
rect 63982 400 64258 430
rect 64374 400 64650 430
rect 64766 400 65042 430
rect 65158 400 65434 430
rect 65550 400 65826 430
rect 65942 400 66218 430
rect 66334 400 66610 430
rect 66726 400 67002 430
rect 67118 400 67394 430
rect 67510 400 67786 430
rect 67902 400 68178 430
rect 68294 400 68570 430
rect 68686 400 68962 430
rect 69078 400 69354 430
rect 69470 400 69746 430
rect 69862 400 70138 430
rect 70254 400 70530 430
rect 70646 400 70922 430
rect 71038 400 71314 430
rect 71430 400 71706 430
rect 71822 400 72098 430
rect 72214 400 72490 430
rect 72606 400 72882 430
rect 72998 400 73274 430
rect 73390 400 73666 430
rect 73782 400 74058 430
rect 74174 400 74450 430
rect 74566 400 74842 430
rect 74958 400 75234 430
rect 75350 400 75626 430
rect 75742 400 76018 430
rect 76134 400 76410 430
rect 76526 400 76802 430
rect 76918 400 77194 430
rect 77310 400 77586 430
rect 77702 400 77978 430
rect 78094 400 78370 430
rect 78486 400 78762 430
rect 78878 400 79154 430
rect 79270 400 79546 430
rect 79662 400 79938 430
rect 80054 400 80330 430
rect 80446 400 80722 430
rect 80838 400 81114 430
rect 81230 400 81506 430
rect 81622 400 81898 430
rect 82014 400 82290 430
rect 82406 400 82682 430
rect 82798 400 83074 430
rect 83190 400 83466 430
rect 83582 400 83858 430
rect 83974 400 84250 430
rect 84366 400 84642 430
rect 84758 400 85034 430
rect 85150 400 85426 430
rect 85542 400 85818 430
rect 85934 400 86210 430
rect 86326 400 86602 430
rect 86718 400 86994 430
rect 87110 400 87386 430
rect 87502 400 87778 430
rect 87894 400 88170 430
rect 88286 400 88562 430
rect 88678 400 88954 430
rect 89070 400 89346 430
rect 89462 400 89738 430
rect 89854 400 90130 430
rect 90246 400 90522 430
rect 90638 400 90914 430
rect 91030 400 91306 430
rect 91422 400 91698 430
rect 91814 400 92090 430
rect 92206 400 92482 430
rect 92598 400 92874 430
rect 92990 400 93266 430
rect 93382 400 93658 430
rect 93774 400 94050 430
rect 94166 400 94442 430
rect 94558 400 94834 430
rect 94950 400 95226 430
rect 95342 400 95618 430
rect 95734 400 96010 430
rect 96126 400 96402 430
rect 96518 400 96794 430
rect 96910 400 97186 430
rect 97302 400 97578 430
rect 97694 400 97970 430
rect 98086 400 98362 430
rect 98478 400 98754 430
rect 98870 400 99146 430
rect 99262 400 99538 430
rect 99654 400 99930 430
rect 100046 400 100322 430
rect 100438 400 100714 430
rect 100830 400 101106 430
rect 101222 400 101498 430
rect 101614 400 101890 430
rect 102006 400 102282 430
rect 102398 400 102674 430
rect 102790 400 103066 430
rect 103182 400 103458 430
rect 103574 400 103850 430
rect 103966 400 104242 430
rect 104358 400 104634 430
rect 104750 400 105026 430
rect 105142 400 105418 430
rect 105534 400 105810 430
rect 105926 400 106202 430
rect 106318 400 106594 430
rect 106710 400 106986 430
rect 107102 400 107378 430
rect 107494 400 107770 430
rect 107886 400 108162 430
rect 108278 400 108554 430
rect 108670 400 108946 430
rect 109062 400 109338 430
rect 109454 400 109730 430
rect 109846 400 110122 430
rect 110238 400 110514 430
rect 110630 400 110906 430
rect 111022 400 111298 430
rect 111414 400 111690 430
rect 111806 400 112082 430
rect 112198 400 112474 430
rect 112590 400 112866 430
rect 112982 400 113258 430
rect 113374 400 113650 430
rect 113766 400 114042 430
rect 114158 400 114434 430
rect 114550 400 114826 430
rect 114942 400 115218 430
rect 115334 400 115610 430
rect 115726 400 116002 430
rect 116118 400 116394 430
rect 116510 400 116786 430
rect 116902 400 117178 430
rect 117294 400 117570 430
rect 117686 400 117962 430
rect 118078 400 118354 430
rect 118470 400 118746 430
rect 118862 400 119138 430
rect 119254 400 119530 430
rect 119646 400 119922 430
rect 120038 400 120314 430
rect 120430 400 120706 430
rect 120822 400 121098 430
rect 121214 400 121490 430
rect 121606 400 121882 430
rect 121998 400 122274 430
rect 122390 400 122666 430
rect 122782 400 123058 430
rect 123174 400 123450 430
rect 123566 400 123842 430
rect 123958 400 124234 430
rect 124350 400 124626 430
rect 124742 400 125018 430
rect 125134 400 125410 430
rect 125526 400 125802 430
rect 125918 400 126194 430
rect 126310 400 126586 430
rect 126702 400 126978 430
rect 127094 400 127370 430
rect 127486 400 127762 430
rect 127878 400 128154 430
rect 128270 400 128546 430
rect 128662 400 128938 430
rect 129054 400 129330 430
rect 129446 400 129722 430
rect 129838 400 130114 430
rect 130230 400 130506 430
rect 130622 400 130898 430
rect 131014 400 131290 430
rect 131406 400 131682 430
rect 131798 400 132074 430
rect 132190 400 132466 430
rect 132582 400 132858 430
rect 132974 400 133250 430
rect 133366 400 133642 430
rect 133758 400 134034 430
rect 134150 400 134426 430
rect 134542 400 134818 430
rect 134934 400 135210 430
rect 135326 400 135602 430
rect 135718 400 135994 430
rect 136110 400 136386 430
rect 136502 400 136778 430
rect 136894 400 137170 430
rect 137286 400 137562 430
rect 137678 400 137954 430
rect 138070 400 138346 430
rect 138462 400 138738 430
rect 138854 400 139130 430
rect 139246 400 139522 430
rect 139638 400 139914 430
rect 140030 400 140306 430
rect 140422 400 140698 430
rect 140814 400 141090 430
rect 141206 400 141482 430
rect 141598 400 141874 430
rect 141990 400 142266 430
rect 142382 400 142658 430
rect 142774 400 143050 430
rect 143166 400 143442 430
rect 143558 400 143834 430
rect 143950 400 144226 430
rect 144342 400 144618 430
rect 144734 400 145010 430
rect 145126 400 145402 430
rect 145518 400 145794 430
rect 145910 400 146186 430
rect 146302 400 146578 430
rect 146694 400 146970 430
rect 147086 400 147362 430
rect 147478 400 147754 430
rect 147870 400 148146 430
rect 148262 400 148538 430
rect 148654 400 148930 430
rect 149046 400 149322 430
rect 149438 400 149714 430
rect 149830 400 150106 430
rect 150222 400 150498 430
rect 150614 400 150890 430
rect 151006 400 151282 430
rect 151398 400 151674 430
rect 151790 400 152066 430
rect 152182 400 152458 430
rect 152574 400 152850 430
rect 152966 400 153242 430
rect 153358 400 153634 430
rect 153750 400 154026 430
rect 154142 400 154418 430
rect 154534 400 154810 430
rect 154926 400 155202 430
rect 155318 400 155594 430
rect 155710 400 155986 430
rect 156102 400 156378 430
rect 156494 400 156770 430
rect 156886 400 157162 430
rect 157278 400 157554 430
rect 157670 400 157946 430
rect 158062 400 158338 430
rect 158454 400 158730 430
rect 158846 400 159122 430
rect 159238 400 159514 430
rect 159630 400 159906 430
rect 160022 400 160298 430
rect 160414 400 160690 430
rect 160806 400 161082 430
rect 161198 400 161474 430
rect 161590 400 161866 430
rect 161982 400 162258 430
rect 162374 400 162650 430
rect 162766 400 163042 430
rect 163158 400 163434 430
rect 163550 400 163826 430
rect 163942 400 164218 430
rect 164334 400 164610 430
rect 164726 400 165002 430
rect 165118 400 165394 430
rect 165510 400 165786 430
rect 165902 400 166178 430
rect 166294 400 166570 430
rect 166686 400 166962 430
rect 167078 400 167354 430
rect 167470 400 167746 430
rect 167862 400 168138 430
rect 168254 400 168530 430
rect 168646 400 168922 430
rect 169038 400 169314 430
rect 169430 400 169706 430
rect 169822 400 170098 430
rect 170214 400 170490 430
rect 170606 400 170882 430
rect 170998 400 171274 430
rect 171390 400 171666 430
rect 171782 400 172058 430
rect 172174 400 172450 430
rect 172566 400 172842 430
rect 172958 400 173234 430
rect 173350 400 173626 430
rect 173742 400 174018 430
rect 174134 400 174410 430
rect 174526 400 174802 430
rect 174918 400 175194 430
rect 175310 400 175586 430
rect 175702 400 175978 430
rect 176094 400 176370 430
rect 176486 400 176762 430
rect 176878 400 177154 430
rect 177270 400 177546 430
rect 177662 400 177938 430
rect 178054 400 178330 430
rect 178446 400 178722 430
rect 178838 400 179114 430
rect 179230 400 179506 430
rect 179622 400 179898 430
rect 180014 400 180290 430
rect 180406 400 180682 430
rect 180798 400 181074 430
rect 181190 400 181466 430
rect 181582 400 181858 430
rect 181974 400 182250 430
rect 182366 400 182642 430
rect 182758 400 183034 430
rect 183150 400 183426 430
rect 183542 400 183818 430
rect 183934 400 184210 430
rect 184326 400 184602 430
rect 184718 400 184994 430
rect 185110 400 185386 430
rect 185502 400 185778 430
rect 185894 400 186170 430
rect 186286 400 186562 430
rect 186678 400 186954 430
rect 187070 400 187346 430
rect 187462 400 187738 430
rect 187854 400 188130 430
rect 188246 400 188522 430
rect 188638 400 188914 430
rect 189030 400 189306 430
rect 189422 400 189698 430
rect 189814 400 190090 430
rect 190206 400 190482 430
rect 190598 400 190874 430
rect 190990 400 191266 430
rect 191382 400 191658 430
rect 191774 400 192050 430
rect 192166 400 192442 430
rect 192558 400 192834 430
rect 192950 400 193226 430
rect 193342 400 193618 430
rect 193734 400 194010 430
rect 194126 400 194402 430
rect 194518 400 194794 430
rect 194910 400 195186 430
rect 195302 400 195578 430
rect 195694 400 195970 430
rect 196086 400 196362 430
rect 196478 400 198170 430
<< obsm3 >>
rect 2233 1554 196943 148190
<< metal4 >>
rect 2224 1538 2384 148206
rect 9904 1538 10064 148206
rect 17584 1538 17744 148206
rect 25264 1538 25424 148206
rect 32944 1538 33104 148206
rect 40624 1538 40784 148206
rect 48304 1538 48464 148206
rect 55984 1538 56144 148206
rect 63664 1538 63824 148206
rect 71344 1538 71504 148206
rect 79024 1538 79184 148206
rect 86704 1538 86864 148206
rect 94384 1538 94544 148206
rect 102064 1538 102224 148206
rect 109744 1538 109904 148206
rect 117424 1538 117584 148206
rect 125104 1538 125264 148206
rect 132784 1538 132944 148206
rect 140464 1538 140624 148206
rect 148144 1538 148304 148206
rect 155824 1538 155984 148206
rect 163504 1538 163664 148206
rect 171184 1538 171344 148206
rect 178864 1538 179024 148206
rect 186544 1538 186704 148206
rect 194224 1538 194384 148206
<< obsm4 >>
rect 47054 105849 48274 141279
rect 48494 105849 55954 141279
rect 56174 105849 63634 141279
rect 63854 105849 71314 141279
rect 71534 105849 78994 141279
rect 79214 105849 86674 141279
rect 86894 105849 94354 141279
rect 94574 105849 102034 141279
rect 102254 105849 109714 141279
rect 109934 105849 117394 141279
rect 117614 105849 125074 141279
rect 125294 105849 131866 141279
<< labels >>
rlabel metal2 s 1848 149600 1904 150000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 53928 149600 53984 150000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 59136 149600 59192 150000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 64344 149600 64400 150000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 69552 149600 69608 150000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 74760 149600 74816 150000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 79968 149600 80024 150000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 85176 149600 85232 150000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 90384 149600 90440 150000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 95592 149600 95648 150000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 100800 149600 100856 150000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 7056 149600 7112 150000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 106008 149600 106064 150000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 111216 149600 111272 150000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 116424 149600 116480 150000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 121632 149600 121688 150000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 126840 149600 126896 150000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 132048 149600 132104 150000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 137256 149600 137312 150000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 142464 149600 142520 150000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 147672 149600 147728 150000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 152880 149600 152936 150000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 12264 149600 12320 150000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 158088 149600 158144 150000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 163296 149600 163352 150000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 168504 149600 168560 150000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 173712 149600 173768 150000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 178920 149600 178976 150000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 184128 149600 184184 150000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 189336 149600 189392 150000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 194544 149600 194600 150000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 17472 149600 17528 150000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 22680 149600 22736 150000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 27888 149600 27944 150000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 33096 149600 33152 150000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 38304 149600 38360 150000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 43512 149600 43568 150000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 48720 149600 48776 150000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3584 149600 3640 150000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 55664 149600 55720 150000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 60872 149600 60928 150000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 66080 149600 66136 150000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 71288 149600 71344 150000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 76496 149600 76552 150000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 81704 149600 81760 150000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 86912 149600 86968 150000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 92120 149600 92176 150000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 97328 149600 97384 150000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 102536 149600 102592 150000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 8792 149600 8848 150000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 107744 149600 107800 150000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 112952 149600 113008 150000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 118160 149600 118216 150000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 123368 149600 123424 150000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 128576 149600 128632 150000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 133784 149600 133840 150000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 138992 149600 139048 150000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 144200 149600 144256 150000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 149408 149600 149464 150000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 154616 149600 154672 150000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 14000 149600 14056 150000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 159824 149600 159880 150000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 165032 149600 165088 150000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 170240 149600 170296 150000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 175448 149600 175504 150000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 180656 149600 180712 150000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 185864 149600 185920 150000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 191072 149600 191128 150000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 196280 149600 196336 150000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 19208 149600 19264 150000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 24416 149600 24472 150000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 29624 149600 29680 150000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 34832 149600 34888 150000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 40040 149600 40096 150000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 45248 149600 45304 150000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 50456 149600 50512 150000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 5320 149600 5376 150000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 57400 149600 57456 150000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 62608 149600 62664 150000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 67816 149600 67872 150000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 73024 149600 73080 150000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 78232 149600 78288 150000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 83440 149600 83496 150000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 88648 149600 88704 150000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 93856 149600 93912 150000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 99064 149600 99120 150000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 104272 149600 104328 150000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 10528 149600 10584 150000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 109480 149600 109536 150000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 114688 149600 114744 150000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 119896 149600 119952 150000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 125104 149600 125160 150000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 130312 149600 130368 150000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 135520 149600 135576 150000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 140728 149600 140784 150000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 145936 149600 145992 150000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 151144 149600 151200 150000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 156352 149600 156408 150000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 15736 149600 15792 150000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 161560 149600 161616 150000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 166768 149600 166824 150000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 171976 149600 172032 150000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 177184 149600 177240 150000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 182392 149600 182448 150000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 187600 149600 187656 150000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 192808 149600 192864 150000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 198016 149600 198072 150000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 20944 149600 21000 150000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 26152 149600 26208 150000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 31360 149600 31416 150000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 36568 149600 36624 150000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 41776 149600 41832 150000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 46984 149600 47040 150000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 52192 149600 52248 150000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 195608 0 195664 400 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 196000 0 196056 400 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 196392 0 196448 400 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 45080 0 45136 400 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 162680 0 162736 400 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 163856 0 163912 400 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 165032 0 165088 400 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 166208 0 166264 400 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 167384 0 167440 400 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 168560 0 168616 400 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 169736 0 169792 400 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 170912 0 170968 400 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 172088 0 172144 400 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 173264 0 173320 400 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 56840 0 56896 400 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 174440 0 174496 400 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 175616 0 175672 400 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 176792 0 176848 400 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 177968 0 178024 400 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 179144 0 179200 400 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 180320 0 180376 400 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 181496 0 181552 400 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 182672 0 182728 400 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 183848 0 183904 400 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 185024 0 185080 400 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 58016 0 58072 400 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 186200 0 186256 400 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 187376 0 187432 400 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 188552 0 188608 400 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 189728 0 189784 400 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 190904 0 190960 400 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 192080 0 192136 400 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 193256 0 193312 400 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 194432 0 194488 400 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 59192 0 59248 400 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 60368 0 60424 400 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 61544 0 61600 400 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 62720 0 62776 400 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 63896 0 63952 400 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 65072 0 65128 400 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 66248 0 66304 400 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 67424 0 67480 400 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 46256 0 46312 400 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 68600 0 68656 400 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 69776 0 69832 400 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 70952 0 71008 400 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 72128 0 72184 400 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 73304 0 73360 400 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 74480 0 74536 400 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 75656 0 75712 400 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 76832 0 76888 400 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 78008 0 78064 400 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 79184 0 79240 400 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 47432 0 47488 400 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 80360 0 80416 400 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 81536 0 81592 400 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 82712 0 82768 400 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 83888 0 83944 400 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 85064 0 85120 400 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 86240 0 86296 400 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 87416 0 87472 400 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 88592 0 88648 400 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 89768 0 89824 400 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 90944 0 91000 400 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 48608 0 48664 400 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 92120 0 92176 400 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 93296 0 93352 400 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 94472 0 94528 400 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 95648 0 95704 400 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 96824 0 96880 400 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 98000 0 98056 400 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 99176 0 99232 400 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 100352 0 100408 400 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 101528 0 101584 400 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 102704 0 102760 400 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 49784 0 49840 400 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 103880 0 103936 400 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 105056 0 105112 400 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 106232 0 106288 400 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 107408 0 107464 400 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 108584 0 108640 400 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 109760 0 109816 400 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 110936 0 110992 400 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 112112 0 112168 400 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 113288 0 113344 400 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 114464 0 114520 400 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 50960 0 51016 400 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 115640 0 115696 400 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 116816 0 116872 400 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 117992 0 118048 400 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 119168 0 119224 400 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 120344 0 120400 400 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 121520 0 121576 400 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 122696 0 122752 400 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 123872 0 123928 400 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 125048 0 125104 400 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 126224 0 126280 400 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 52136 0 52192 400 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 127400 0 127456 400 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 128576 0 128632 400 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 129752 0 129808 400 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 130928 0 130984 400 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 132104 0 132160 400 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 133280 0 133336 400 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 134456 0 134512 400 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 135632 0 135688 400 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 136808 0 136864 400 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 137984 0 138040 400 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 53312 0 53368 400 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 139160 0 139216 400 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 140336 0 140392 400 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 141512 0 141568 400 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 142688 0 142744 400 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 143864 0 143920 400 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 145040 0 145096 400 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 146216 0 146272 400 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 147392 0 147448 400 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 148568 0 148624 400 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 149744 0 149800 400 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 54488 0 54544 400 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 150920 0 150976 400 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 152096 0 152152 400 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 153272 0 153328 400 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 154448 0 154504 400 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 155624 0 155680 400 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 156800 0 156856 400 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 157976 0 158032 400 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 159152 0 159208 400 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 160328 0 160384 400 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 161504 0 161560 400 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 55664 0 55720 400 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 45472 0 45528 400 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 163072 0 163128 400 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 164248 0 164304 400 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 165424 0 165480 400 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 166600 0 166656 400 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 167776 0 167832 400 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 168952 0 169008 400 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 170128 0 170184 400 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 171304 0 171360 400 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 172480 0 172536 400 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 173656 0 173712 400 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 57232 0 57288 400 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 174832 0 174888 400 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 176008 0 176064 400 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 177184 0 177240 400 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 178360 0 178416 400 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 179536 0 179592 400 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 180712 0 180768 400 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 181888 0 181944 400 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 183064 0 183120 400 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 184240 0 184296 400 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 185416 0 185472 400 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 58408 0 58464 400 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 186592 0 186648 400 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 187768 0 187824 400 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 188944 0 189000 400 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 190120 0 190176 400 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 191296 0 191352 400 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 192472 0 192528 400 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 193648 0 193704 400 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 194824 0 194880 400 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 59584 0 59640 400 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 60760 0 60816 400 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 61936 0 61992 400 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 63112 0 63168 400 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 64288 0 64344 400 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 65464 0 65520 400 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 66640 0 66696 400 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 67816 0 67872 400 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 46648 0 46704 400 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 68992 0 69048 400 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 70168 0 70224 400 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 71344 0 71400 400 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 72520 0 72576 400 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 73696 0 73752 400 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 74872 0 74928 400 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 76048 0 76104 400 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 77224 0 77280 400 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 78400 0 78456 400 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 79576 0 79632 400 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 47824 0 47880 400 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 80752 0 80808 400 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 81928 0 81984 400 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 83104 0 83160 400 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 84280 0 84336 400 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 85456 0 85512 400 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 86632 0 86688 400 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 87808 0 87864 400 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 88984 0 89040 400 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 90160 0 90216 400 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 91336 0 91392 400 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 49000 0 49056 400 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 92512 0 92568 400 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 93688 0 93744 400 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 94864 0 94920 400 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 96040 0 96096 400 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 97216 0 97272 400 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 98392 0 98448 400 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 99568 0 99624 400 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 100744 0 100800 400 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 101920 0 101976 400 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 103096 0 103152 400 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 50176 0 50232 400 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 104272 0 104328 400 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 105448 0 105504 400 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 106624 0 106680 400 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 107800 0 107856 400 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 108976 0 109032 400 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 110152 0 110208 400 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 111328 0 111384 400 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 112504 0 112560 400 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 113680 0 113736 400 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 114856 0 114912 400 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 51352 0 51408 400 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 116032 0 116088 400 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 117208 0 117264 400 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 118384 0 118440 400 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 119560 0 119616 400 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 120736 0 120792 400 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 121912 0 121968 400 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 123088 0 123144 400 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 124264 0 124320 400 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 125440 0 125496 400 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 126616 0 126672 400 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 52528 0 52584 400 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 127792 0 127848 400 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 128968 0 129024 400 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 130144 0 130200 400 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 131320 0 131376 400 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 132496 0 132552 400 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 133672 0 133728 400 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 134848 0 134904 400 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 136024 0 136080 400 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 137200 0 137256 400 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 138376 0 138432 400 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 53704 0 53760 400 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 139552 0 139608 400 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 140728 0 140784 400 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 141904 0 141960 400 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 143080 0 143136 400 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 144256 0 144312 400 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 145432 0 145488 400 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 146608 0 146664 400 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 147784 0 147840 400 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 148960 0 149016 400 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 150136 0 150192 400 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 54880 0 54936 400 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 151312 0 151368 400 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 152488 0 152544 400 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 153664 0 153720 400 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 154840 0 154896 400 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 156016 0 156072 400 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 157192 0 157248 400 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 158368 0 158424 400 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 159544 0 159600 400 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 160720 0 160776 400 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 161896 0 161952 400 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 56056 0 56112 400 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 45864 0 45920 400 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 163464 0 163520 400 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 164640 0 164696 400 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 165816 0 165872 400 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 166992 0 167048 400 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 168168 0 168224 400 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 169344 0 169400 400 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 170520 0 170576 400 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 171696 0 171752 400 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 172872 0 172928 400 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 174048 0 174104 400 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 57624 0 57680 400 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 175224 0 175280 400 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 176400 0 176456 400 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 177576 0 177632 400 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 178752 0 178808 400 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 179928 0 179984 400 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 181104 0 181160 400 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 182280 0 182336 400 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 183456 0 183512 400 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 184632 0 184688 400 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 185808 0 185864 400 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 58800 0 58856 400 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 186984 0 187040 400 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 188160 0 188216 400 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 189336 0 189392 400 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 190512 0 190568 400 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 191688 0 191744 400 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 192864 0 192920 400 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 194040 0 194096 400 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 195216 0 195272 400 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 59976 0 60032 400 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 61152 0 61208 400 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 62328 0 62384 400 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 63504 0 63560 400 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 64680 0 64736 400 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 65856 0 65912 400 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 67032 0 67088 400 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 68208 0 68264 400 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 47040 0 47096 400 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 69384 0 69440 400 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 70560 0 70616 400 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 71736 0 71792 400 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 72912 0 72968 400 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 74088 0 74144 400 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 75264 0 75320 400 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 76440 0 76496 400 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 77616 0 77672 400 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 78792 0 78848 400 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 79968 0 80024 400 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 48216 0 48272 400 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 81144 0 81200 400 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 82320 0 82376 400 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 83496 0 83552 400 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 84672 0 84728 400 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 85848 0 85904 400 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 87024 0 87080 400 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 88200 0 88256 400 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 89376 0 89432 400 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 90552 0 90608 400 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 91728 0 91784 400 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 49392 0 49448 400 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 92904 0 92960 400 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 94080 0 94136 400 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 95256 0 95312 400 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 96432 0 96488 400 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 97608 0 97664 400 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 98784 0 98840 400 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 99960 0 100016 400 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 101136 0 101192 400 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 102312 0 102368 400 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 103488 0 103544 400 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 50568 0 50624 400 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 104664 0 104720 400 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 105840 0 105896 400 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 107016 0 107072 400 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 108192 0 108248 400 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 109368 0 109424 400 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 110544 0 110600 400 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 111720 0 111776 400 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 112896 0 112952 400 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 114072 0 114128 400 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 115248 0 115304 400 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 51744 0 51800 400 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 116424 0 116480 400 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 117600 0 117656 400 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 118776 0 118832 400 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 119952 0 120008 400 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 121128 0 121184 400 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 122304 0 122360 400 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 123480 0 123536 400 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 124656 0 124712 400 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 125832 0 125888 400 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 127008 0 127064 400 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 52920 0 52976 400 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 128184 0 128240 400 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 129360 0 129416 400 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 130536 0 130592 400 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 131712 0 131768 400 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 132888 0 132944 400 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 134064 0 134120 400 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 135240 0 135296 400 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 136416 0 136472 400 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 137592 0 137648 400 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 138768 0 138824 400 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 54096 0 54152 400 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 139944 0 140000 400 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 141120 0 141176 400 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 142296 0 142352 400 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 143472 0 143528 400 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 144648 0 144704 400 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 145824 0 145880 400 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 147000 0 147056 400 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 148176 0 148232 400 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 149352 0 149408 400 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 150528 0 150584 400 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 55272 0 55328 400 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 151704 0 151760 400 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 152880 0 152936 400 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 154056 0 154112 400 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 155232 0 155288 400 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 156408 0 156464 400 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 157584 0 157640 400 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 158760 0 158816 400 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 159936 0 159992 400 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 161112 0 161168 400 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 162288 0 162344 400 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 56448 0 56504 400 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 2224 1538 2384 148206 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 148206 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 148206 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 148206 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 148206 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 148206 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 148206 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 148206 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 148206 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 148206 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 148206 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 148206 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 148206 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 148206 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 148206 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 148206 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 148206 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 148206 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 148206 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 148206 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 148206 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 148206 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 148206 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 148206 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 148206 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 194224 1538 194384 148206 6 vssd1
port 503 nsew ground bidirectional
rlabel metal2 s 3528 0 3584 400 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 3920 0 3976 400 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 4312 0 4368 400 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 5880 0 5936 400 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 19208 0 19264 400 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 20384 0 20440 400 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 21560 0 21616 400 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 22736 0 22792 400 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 23912 0 23968 400 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 25088 0 25144 400 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 26264 0 26320 400 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 27440 0 27496 400 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 28616 0 28672 400 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 29792 0 29848 400 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 7448 0 7504 400 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 30968 0 31024 400 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 32144 0 32200 400 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 33320 0 33376 400 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 34496 0 34552 400 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 35672 0 35728 400 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 36848 0 36904 400 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 38024 0 38080 400 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 39200 0 39256 400 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 40376 0 40432 400 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 41552 0 41608 400 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 9016 0 9072 400 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 42728 0 42784 400 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 43904 0 43960 400 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 10584 0 10640 400 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 12152 0 12208 400 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 13328 0 13384 400 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 14504 0 14560 400 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 15680 0 15736 400 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 16856 0 16912 400 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 18032 0 18088 400 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 4704 0 4760 400 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 6272 0 6328 400 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 19600 0 19656 400 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 20776 0 20832 400 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 21952 0 22008 400 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 23128 0 23184 400 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 24304 0 24360 400 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 25480 0 25536 400 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 26656 0 26712 400 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 27832 0 27888 400 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 29008 0 29064 400 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 30184 0 30240 400 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 7840 0 7896 400 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 31360 0 31416 400 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 32536 0 32592 400 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 33712 0 33768 400 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 34888 0 34944 400 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 36064 0 36120 400 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 37240 0 37296 400 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 38416 0 38472 400 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 39592 0 39648 400 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 40768 0 40824 400 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 41944 0 42000 400 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 9408 0 9464 400 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 43120 0 43176 400 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 44296 0 44352 400 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 10976 0 11032 400 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 12544 0 12600 400 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 13720 0 13776 400 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 14896 0 14952 400 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 16072 0 16128 400 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 17248 0 17304 400 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 18424 0 18480 400 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 6664 0 6720 400 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 19992 0 20048 400 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 21168 0 21224 400 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 22344 0 22400 400 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 23520 0 23576 400 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 24696 0 24752 400 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 25872 0 25928 400 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 27048 0 27104 400 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 28224 0 28280 400 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 29400 0 29456 400 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 30576 0 30632 400 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 8232 0 8288 400 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 31752 0 31808 400 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 32928 0 32984 400 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 34104 0 34160 400 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 35280 0 35336 400 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 36456 0 36512 400 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 37632 0 37688 400 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 38808 0 38864 400 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 39984 0 40040 400 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 41160 0 41216 400 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 42336 0 42392 400 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 9800 0 9856 400 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 43512 0 43568 400 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 44688 0 44744 400 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 11368 0 11424 400 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 12936 0 12992 400 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 14112 0 14168 400 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 15288 0 15344 400 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 16464 0 16520 400 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 17640 0 17696 400 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 18816 0 18872 400 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 7056 0 7112 400 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 8624 0 8680 400 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 10192 0 10248 400 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 11760 0 11816 400 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 5096 0 5152 400 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 5488 0 5544 400 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 200000 150000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 17088734
string GDS_FILE /home/radhe/tapeout_projects/radhe_gf180nm/openlane/user_proj_example/runs/22_12_05_06_53/results/signoff/user_proj_example.magic.gds
string GDS_START 285444
<< end >>

