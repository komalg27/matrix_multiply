* NGSPICE file created from matrix_multiply.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_20 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_20 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

.subckt matrix_multiply clk execute input_val[0] input_val[1] input_val[2] input_val[3]
+ input_val[4] input_val[5] input_val[6] input_val[7] reset result[0] result[10] result[11]
+ result[12] result[13] result[14] result[15] result[16] result[1] result[2] result[3]
+ result[4] result[5] result[6] result[7] result[8] result[9] sel_in[0] sel_in[1]
+ sel_in[2] sel_out[0] sel_out[1] vccd1 vssd1
XFILLER_140_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5417__B1 _0712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5968__A1 _1896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4640__A1 _3181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6845_ _0028_ net11 net1 A\[3\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6776_ _2673_ _2200_ _2724_ _2729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5196__A2 _1054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6393__A1 _2361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3988_ _0784_ _3079_ _3140_ _3148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_5727_ _1336_ _1343_ _1639_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_136_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6160__I _1482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5658_ _1505_ _1562_ _1563_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4609_ _0397_ _0398_ _0433_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5589_ _1486_ _0998_ _1437_ _0999_ _1487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_123_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6448__A2 _2427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4459__A1 _2930_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5423__A3 _1285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6860__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5187__A2 _1044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4934__A2 _0766_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4698__A1 _3371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3673__A2 _2832_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6611__A2 _1187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4960_ _0748_ _0752_ _0794_ _0796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4622__A1 _0315_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3911_ _0718_ _2939_ _3071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4891_ _0714_ _0719_ _0720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6851__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3976__A3 _3135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6630_ _1661_ _1804_ _1586_ _2617_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3842_ _3000_ _3001_ _3002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5178__A2 _0941_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6561_ _1749_ _1759_ _2547_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3773_ _2932_ _2933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4925__A2 _0755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5512_ _1401_ _1363_ _1402_ _1376_ _1403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6127__A1 _1562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6492_ _2275_ _2474_ _2475_ _2264_ _2476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_121_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5443_ _1281_ _1326_ _1327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5350__A2 _1223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5374_ _1250_ _1248_ _3270_ _3272_ _1251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_99_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4325_ _3382_ _0149_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4256_ _0079_ _0080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5102__A2 _0951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4310__B1 _2988_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4187_ _3346_ _2786_ _3347_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3779__I _1081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6602__A2 _2581_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4613__A1 _0424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6842__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5169__A2 _0931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6828_ _0011_ net11 net1 A\[1\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6759_ _2654_ _2703_ _2717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6669__A2 _2632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3655__A2 _2813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6833__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4907__A2 _0736_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3591__A1 _2179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3894__A2 _3052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4110_ _3269_ _3270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5090_ _0935_ _0936_ _0939_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_111_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5096__A1 _0868_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4041_ _3199_ _3200_ _3201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_110_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5992_ _3220_ _3287_ _1930_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_91_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4943_ _0775_ _0776_ _0777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6824__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4874_ _0683_ _0698_ _0700_ _0701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_32_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6613_ _2597_ _2598_ _2599_ _2491_ _2264_ _2600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3825_ _2984_ _2985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4223__I _3382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6544_ _3180_ _3191_ _2529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_118_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3756_ _2858_ _2871_ _2915_ _2916_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6475_ _2199_ _2202_ _2458_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3687_ _2842_ _2846_ _2847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_134_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5426_ _0072_ _0684_ _1308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4126__A3 _3285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6520__A1 _2368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5357_ _0834_ _1231_ _1232_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_102_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4308_ _3350_ _2863_ _0132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5288_ _1062_ _1156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4239_ A\[0\]\[2\] _3399_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3637__A2 _1554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4062__A2 _3221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6339__A1 _2306_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5011__A1 _0847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6817__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5562__A2 _0473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3573__A1 _2376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5314__A2 _1120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6511__A1 _2421_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4668__A4 _0472_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3876__A2 _3032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3628__A2 _0861_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6724__S _2692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6578__A1 _1794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4589__B1 _0354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3800__A2 _2704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3610_ _2768_ _2769_ _2770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4590_ _0410_ _0412_ _0413_ _0404_ _0414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_128_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3564__A1 _2408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3541_ _2179_ _1960_ _2212_ _2223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_116_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6260_ _2188_ _1922_ _2222_ _2224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5305__A2 _1135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3472_ _0861_ _0993_ _1466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5211_ _1009_ _3108_ _1072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5856__A3 _1780_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6191_ _1940_ _1973_ _2148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3867__A2 _3026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5142_ _0975_ _0995_ _0996_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_111_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5069__A1 _0682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5073_ _0694_ _3044_ _3271_ _0917_ _0920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4816__A1 _0631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4024_ _3182_ _1829_ _3183_ _3184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_49_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6569__A1 _3199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5975_ _1909_ _1910_ _1911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4926_ _0678_ _0756_ _0757_ _0758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4857_ _0681_ _0682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3808_ _2879_ _2967_ _2430_ _2812_ _2968_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4788_ B\[0\]\[6\] _0612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4888__I B\[0\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6527_ _3076_ _3187_ _2512_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3739_ _2875_ _2898_ _2899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_118_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6458_ _2379_ _2384_ _2439_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5409_ _0731_ _0327_ _1289_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6809__S _2751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6389_ _2229_ _2362_ _2363_ _2364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3858__A2 _0784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5480__A1 _1362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4128__I net16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4035__A2 _3179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5783__A2 _1699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3794__A1 _2941_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5535__A2 _0088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4743__B1 _2813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5299__A1 _1124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3849__A2 _2961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6263__A3 _2222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5471__A1 _0649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3877__I _2398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5223__A1 _0973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5760_ _1672_ _1674_ _1676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4711_ _1785_ _0420_ _0535_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5691_ _1599_ _1600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4642_ _0464_ _0465_ _0466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3537__A1 _2157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4573_ _0393_ _0394_ _0396_ _0384_ _0397_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_7_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6312_ _2279_ _2066_ _2280_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4501__I _0133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3524_ B\[1\]\[2\] _2037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6243_ _2197_ _2204_ _2205_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3455_ _1257_ _1268_ _1279_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6174_ _2061_ _2128_ _2129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_97_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5125_ _0875_ _0882_ _0977_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_131_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5056_ _0899_ _0900_ _0901_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4265__A2 _3033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4007_ _3161_ _3162_ _3157_ _3167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_84_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4392__B _0215_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4017__A2 _3172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6163__I _2115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5958_ _1885_ _1891_ _1892_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_90_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5765__A2 _0420_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3776__A1 _2934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4909_ _0714_ _0719_ _0739_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5889_ _0420_ _1817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3700__A1 _1444_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5453__A1 _1310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5205__A1 _1064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5508__A2 _1397_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4192__A1 _3351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5692__A1 _1597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5152__I _0800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4247__A2 _0070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5444__A1 _0623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4991__I _0829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5995__A2 _3286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6861_ _0044_ net11 net1 B\[1\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5812_ _1729_ _1732_ _1733_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3400__I net15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6792_ _1595_ _2645_ _2738_ _2741_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5743_ _1655_ _1656_ _1657_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6711__I _2685_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5674_ _1534_ _1571_ _1580_ _1581_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_30_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4625_ _0436_ _0447_ _0448_ _0449_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5327__I _0668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4556_ _0377_ _0378_ _0380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3507_ _1774_ _1840_ _1851_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_1_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4487_ _3344_ _0305_ _3312_ _0311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_143_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6226_ _2183_ _2185_ _2186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_3438_ _1070_ _1081_ _1092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5683__A1 _0307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6157_ _2064_ _2072_ _2110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5108_ _0837_ _0958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6088_ _1195_ _2033_ _2034_ _2035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5435__A1 _1314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5039_ _0880_ _0881_ _0882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_39_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput20 net20 result[12] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput31 net31 result[7] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_134_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6710__I1 _3247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5426__A1 _0072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5977__A2 _2908_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3988__A1 _0784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5729__A2 _1639_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4410_ _0217_ _0232_ _0233_ _0234_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5390_ _1267_ _1269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5901__A2 _1549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4341_ _0164_ _1938_ _0165_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4986__I _0613_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4272_ _0093_ _0094_ _0092_ _0096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6011_ _1943_ _1950_ _1951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5665__A1 _1553_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4468__A2 _2945_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5417__A1 _0073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6614__B1 _2595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5417__B2 _3380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6706__I _2681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6090__A1 _2027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4640__A2 _0190_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6844_ _0027_ net11 net1 A\[3\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3987_ _3139_ _3146_ _3147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6775_ _2728_ _0046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5726_ _1607_ _1628_ _1636_ _1637_ _1638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_136_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5657_ _0836_ _3334_ _1562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6850__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4156__A1 A\[1\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4608_ _0321_ _0322_ _0432_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5588_ _0075_ _1486_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6597__B _2582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4539_ _0331_ _0352_ _0361_ _0362_ _0363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_105_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4459__A2 _0282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6209_ _2165_ _2166_ _2167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5408__A1 _0635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4136__I _3295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6384__A2 _2257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5592__B1 _0548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5895__A1 _1556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5647__A1 _1545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4870__A2 _0688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3910_ _3068_ _3069_ _3070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4890_ _0711_ _0715_ _0717_ _0719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__3830__B1 _2922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3841_ _2991_ _2992_ _3001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3885__I _2113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6375__A2 _2160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5178__A3 _0907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6873__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6560_ _1267_ _2546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3772_ _2931_ _2932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5511_ _1375_ _1371_ _1402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6491_ _2401_ _2404_ _2475_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6127__A2 _1836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4138__A1 _2942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5442_ A\[0\]\[1\] _0627_ _1326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5373_ _0733_ _1250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5350__A3 _3246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4324_ _0111_ _1191_ _0148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5638__A1 _1539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4255_ A\[0\]\[6\] _0079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4310__A1 _3351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4310__B2 _0133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4186_ _3345_ _3346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6063__A1 _0834_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4613__A2 _0427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6827_ _0010_ net11 net1 A\[1\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4377__A1 _1565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6758_ _2716_ _0039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5709_ _0668_ _0342_ _1619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6689_ _2667_ _0012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4301__A1 _0091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3655__A3 _2814_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4604__A2 _0424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5801__A1 _1717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4368__A1 _2921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3591__A2 _2684_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5868__A1 _1761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5868__B2 _1793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6293__A1 _1985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4040_ _3166_ _3195_ _3194_ _3200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_84_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6045__A1 _1238_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5991_ _0696_ _1928_ _1929_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6596__A2 _3209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4942_ _1499_ B\[2\]\[3\] _0776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4873_ _3263_ _0699_ _0700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4504__I _0327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6612_ _0514_ _0519_ _2599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3824_ A\[3\]\[2\] _2984_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5020__A2 _0860_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6543_ _0487_ _0497_ _2226_ _2528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3755_ _2855_ _2872_ _2915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6474_ _2302_ _2316_ _2457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3686_ _2844_ _2845_ _2846_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5425_ _1304_ _1305_ _1306_ _1307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5335__I _3116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4531__A1 _3101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5356_ _2938_ _0958_ _1231_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4307_ _0127_ _0130_ _0131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5287_ _1154_ _1142_ _1155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5087__A2 _0932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4238_ _3378_ _3396_ _3397_ _3398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6166__I _1223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5070__I _0699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4169_ _3262_ _3328_ _3329_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4598__A1 _0414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5011__A2 _0849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4589__A1 _0411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4589__B2 _3039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5250__A2 _1113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3540_ _2048_ _2201_ _2212_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3471_ _1444_ _0817_ _1455_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5305__A3 _1123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5210_ _1065_ _1067_ _1069_ _1071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_143_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6190_ _2145_ _2147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5141_ _3004_ _0970_ _0995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5072_ _0800_ _3108_ _0919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4023_ _3107_ _3170_ _3158_ _3183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6018__A1 _2946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6569__A2 _2147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6813__I0 _1898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5974_ _0552_ _0554_ _1910_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5241__A2 _1102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4925_ _0724_ _0755_ _0757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4856_ B\[0\]\[1\] _0681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3807_ _2190_ _2967_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4787_ _0593_ _0609_ _0610_ _0611_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6526_ _1718_ _1787_ _1788_ _2511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_119_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3738_ _2886_ _2897_ _2898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_107_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6457_ _2383_ _2438_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3669_ _2387_ B\[1\]\[3\] _2829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5408_ _0635_ _3325_ _1288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6388_ _2259_ _2260_ _2258_ _2363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5339_ _0827_ _0842_ _1212_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_88_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4807__A2 _0621_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6009__A1 _3275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3491__A1 _1433_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6804__I0 _3174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4743__A1 _3393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3546__A2 _1158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4743__B2 _0112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5299__A2 _1135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6496__A1 _2437_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6735__S _2698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5471__A2 A\[1\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6420__A1 _1273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4710_ _0259_ _0298_ _0533_ _0534_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4982__A1 _0783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5690_ _0963_ _0313_ _0314_ _0959_ _1599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4641_ _0409_ _0416_ _0403_ _0465_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_128_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4572_ _2983_ _0395_ _3072_ _3367_ _0396_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6311_ _2114_ _2279_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3523_ _1147_ _2026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6487__A1 _1271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3454_ _1169_ _1202_ _1268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6242_ _2199_ _2203_ _2204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_131_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6709__I _2683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6173_ _2126_ _2127_ _2128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5124_ _3005_ _0970_ _0975_ _0976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_84_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5055_ _0587_ _0592_ _0900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4006_ _3155_ _3165_ _3166_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_38_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3473__A1 _1059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5214__A2 _1073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5957_ _0564_ _1890_ _1891_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4908_ _0726_ _0737_ _0738_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5888_ _1814_ _1580_ _1815_ _1816_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4839_ _0611_ _0661_ _0662_ _0663_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4725__A1 _2930_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6509_ _2342_ _2428_ _2494_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3700__A2 B\[3\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5453__A2 _0088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5205__A2 _2932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3767__A2 _2899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4716__A1 _0280_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4192__A2 _1015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6469__A1 _2448_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5141__A1 _3004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5444__A2 _0327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3455__A1 _1257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6860_ _0043_ net11 net1 B\[1\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_62_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5811_ _1731_ _0351_ _0350_ _1140_ _1732_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_62_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6791_ _2740_ _0052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4955__A1 _0635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5742_ _1459_ _1460_ _1656_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5673_ _1578_ _1579_ _1580_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4707__A1 _2909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4624_ _0439_ _0440_ _0448_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4555_ _0377_ _0378_ _0379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3506_ _1785_ _1829_ _1840_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4486_ _0305_ _0306_ _0308_ _0309_ _0310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_89_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6225_ _2184_ _1980_ _2185_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3437_ B\[3\]\[3\] _1081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5683__A2 _0951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6156_ _2107_ _2108_ _2109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5107_ _0955_ _0956_ _0957_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6087_ _1198_ _1263_ _2034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_73_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5435__A2 _1317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5038_ _0602_ _0603_ _0601_ _0881_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA_input11_I reset vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4946__A1 _0764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4410__A3 _0233_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput21 net21 result[13] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput32 net32 result[8] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_27_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3685__A1 _2780_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5428__I _0716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4340_ A\[0\]\[7\] _0164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4271_ _0092_ _0093_ _0094_ _0095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_140_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6010_ _3266_ _1948_ _1950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_80_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input3_I input_val[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5417__A2 _0699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6090__A2 _2030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4640__A3 _0463_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6843_ _0026_ net11 net1 A\[3\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4928__A1 _0654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6774_ _2647_ _2198_ _2724_ _2728_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3986_ _3141_ _3144_ _3145_ _3146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_22_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5725_ _1634_ _1635_ _1637_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5656_ _1228_ _3353_ _1561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4156__A2 _1510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4607_ _0402_ _0429_ _0430_ _0431_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5587_ _1476_ _1484_ _1485_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_117_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4538_ _0359_ _0360_ _0362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3903__A2 _3060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4469_ _0291_ _0292_ _0293_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5656__A2 _3353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6208_ _3275_ _1947_ _2166_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6139_ _1813_ _1861_ _2091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6081__A2 _1262_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4092__A1 _3251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4919__A1 _0622_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4395__A2 _0217_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5592__A1 _1222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5592__B2 _0613_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5344__A1 _0845_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6541__B1 _2526_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3830__A1 _2985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3840_ _2997_ _2999_ _3000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3771_ _2814_ _2931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5510_ _3350_ _0594_ _1401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6490_ _2401_ _2404_ _2474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4997__I _0833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5441_ _1293_ _1324_ _1325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4138__A2 _3297_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5372_ _1247_ _3270_ _3272_ _1248_ _1249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_126_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5350__A4 _3247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4323_ _0093_ _0146_ _0147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5638__A2 _1540_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4254_ _2037_ _0069_ _0078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6864__D _0047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6717__I _2688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4310__A2 _3307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4185_ A\[1\]\[5\] _3345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6063__A2 _2007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6653__S _2638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6826_ _0009_ net11 net1 A\[1\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6757_ _2673_ _2120_ _2712_ _2716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4377__A2 _3308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3969_ _3128_ _3087_ _3129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5708_ _1614_ _1617_ _1618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_109_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6688_ _2665_ _1817_ _2666_ _2667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5639_ _1538_ _1541_ _1542_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_128_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5877__A2 _1801_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3655__A4 _2288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4147__I _0861_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4604__A3 _0427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5801__A2 _1720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3812__A1 _2966_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4368__A2 _0191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5868__A2 _1781_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5990_ _1922_ _1926_ _1928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6840__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4056__A1 _2904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4941_ _2790_ _0649_ _0775_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3803__A1 _2959_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4872_ _0684_ _0699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6611_ _1183_ _1187_ _2043_ _2598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3823_ _1015_ _2983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5556__A1 _1369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6542_ _1784_ _1792_ _2527_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_3754_ _2851_ _2901_ _2913_ _2914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6473_ _2455_ _2456_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3685_ _2780_ _2782_ _2845_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5859__A2 _1780_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5424_ _1299_ _1303_ _1306_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4531__A2 _0354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5355_ _1229_ _3004_ _1230_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6659__I1 _2642_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4306_ _3360_ _0129_ _0130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_88_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5286_ _1073_ _1141_ _1128_ _1154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4237_ _3389_ _3395_ _3397_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4295__A1 _0087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4168_ A\[0\]\[0\] _3328_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4099_ _2964_ _2973_ _3258_ _3259_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4598__A2 _0415_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5547__A1 _1250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6809_ _0319_ _2642_ _2751_ _2752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6863__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4038__A1 _3194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4589__A2 _3043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6306__B _2061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4210__A1 _2921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3470_ A\[3\]\[5\] _1444_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5140_ _0968_ _0978_ _0994_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6266__A2 _2035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5071_ _0917_ _3044_ _0918_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4022_ _3181_ _3182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6018__A2 _1957_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4029__A1 _3172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6813__I1 _2647_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5973_ _0290_ _0553_ _1909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4924_ _0724_ _0755_ _0756_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_21_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4855_ _0626_ _0629_ _0624_ _0680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_138_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6730__I _2691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3806_ _2829_ _2959_ _2965_ _2889_ _2966_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_119_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4786_ _0605_ _0608_ _0610_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6525_ _2400_ _2510_ net17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3737_ _2888_ _2896_ _2897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_118_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6456_ _2159_ _2161_ _2437_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_118_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3668_ _2824_ _2827_ _2828_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_106_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5407_ _0286_ _0615_ _1287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6387_ _2259_ _2260_ _2258_ _2362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3599_ _2627_ _1169_ _2365_ _2758_ _2759_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_121_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5338_ _0835_ _1210_ _1211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4268__A1 A\[1\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5269_ _1127_ _1133_ _1134_ _1135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6804__I1 _2637_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5768__A1 _3328_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3469__C _1422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4743__A2 _2812_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5759__A1 _0387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6420__A2 _2336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4982__A2 _0804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4640_ _3181_ _0190_ _0463_ _0464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4571_ _0392_ _0395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6310_ _1845_ _2069_ _2123_ _2125_ _2129_ _2278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_3522_ _1982_ _2004_ _2015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6487__A2 _2470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6241_ _2118_ _2198_ _2202_ _2203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3453_ _1235_ _1246_ _1257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6731__I0 _2665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6172_ _1850_ _2068_ _2127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5123_ _0974_ _0975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5054_ _0646_ _0871_ _0899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5998__A1 _1877_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4005_ _3157_ _3163_ _3164_ _3165_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4245__I _3379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5956_ _0568_ _1889_ _1890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_52_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4907_ _0730_ _0736_ _0737_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5887_ _1534_ _1571_ _1815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4838_ _0642_ _0660_ _0662_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_14_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4725__A2 _3245_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4769_ _0587_ _0592_ _0593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_119_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6508_ _2432_ _2493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6439_ _1272_ _2418_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6722__I0 _2652_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5989__A1 _1876_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4661__A1 _0482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4413__A1 _0226_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5913__A1 _1241_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5141__A2 _0970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6746__S _2706_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5810_ _1068_ _1731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_90_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4065__I _2923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6790_ _1596_ _2642_ _2738_ _2740_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5741_ _1624_ _1647_ _1649_ _1651_ _1654_ _1655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__4955__A2 _0734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5672_ _1199_ _0530_ _1579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4623_ _0439_ _0440_ _0447_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5904__A1 _1545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4707__A2 _0530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3409__I B\[3\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4554_ _3372_ _0178_ _0378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3505_ _1818_ _1829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5624__I _1200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4485_ _0189_ _3072_ _0256_ _2983_ _0309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6224_ _1975_ _1978_ _2184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3436_ A\[3\]\[3\] _1070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6656__S _2638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6155_ _2074_ _2086_ _2108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4891__A1 _0714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5106_ _0598_ _0947_ _0877_ _0956_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_111_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6086_ _0945_ _2032_ _2033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_131_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5037_ _0603_ _0876_ _0877_ _0879_ _0880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_100_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6872__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5939_ _0303_ _0524_ _0582_ _1871_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4946__A2 _0779_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6148__A1 _1929_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput22 net22 result[14] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput33 net33 result[9] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_122_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4882__A1 _2704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4634__A1 _0374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6863__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5362__A2 _0860_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4270_ _2763_ A\[0\]\[0\] A\[0\]\[1\] _2762_ _0094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5114__A2 _0964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4873__A1 _3263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3676__A2 _2835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6614__A2 _2592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6854__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6842_ _0025_ net11 net1 A\[3\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6773_ _2727_ _0045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4928__A2 _0658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3985_ _3029_ _3057_ _3145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5050__A1 _0605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5724_ _1634_ _1635_ _1636_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5655_ _0287_ _0830_ _1401_ _1560_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4606_ _0419_ _0428_ _0430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6550__A1 _2268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5586_ _1481_ _1483_ _1484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4537_ _0359_ _0360_ _0361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6302__A1 _2131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4468_ _3346_ _2945_ _2950_ _3351_ _0292_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6207_ _3267_ _1946_ _2165_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3419_ _0872_ _0883_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4399_ _2969_ _2813_ _3323_ _0161_ _0223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6138_ _1816_ _1860_ _2090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5303__B _1172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6605__A2 _1801_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6069_ _1220_ _1234_ _2013_ _2014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6845__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4092__A2 _2949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6369__A1 _1200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4919__A2 _2201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4433__I _0256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5592__A2 _0547_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6541__A1 _2520_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5344__A2 _0862_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4855__A1 _0626_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6309__B _2275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6836__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3830__A2 _2988_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3770_ _1312_ _2930_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5583__A2 _1479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5440_ _1307_ _1322_ _1324_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6532__A1 _2418_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5371_ _0731_ _1248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4322_ _0092_ _0093_ _0094_ _0146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_113_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4253_ _0071_ _0074_ _0076_ _3391_ _0077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_101_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4184_ _3307_ _3313_ _3344_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6827__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6825_ _0008_ net11 net1 A\[1\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__5349__I _1222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6756_ _2715_ _0038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3968_ _3084_ _3085_ _3128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5707_ _1615_ _1616_ _1617_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6687_ _2655_ _2666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_137_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3899_ _3029_ _3057_ _3058_ _3059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6523__A1 _1788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5638_ _1539_ _1540_ _1541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4534__B1 _0357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5569_ _1395_ _1398_ _1465_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3888__A2 _3038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4837__A1 _0642_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6818__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5262__A1 _1065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5317__A2 _1183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4940_ _0771_ _0657_ _0772_ _0774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4871_ _0689_ _2495_ _0698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5005__A1 _0793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6610_ _1183_ _1187_ _2597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3822_ _2786_ _0982_ _2982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3567__A1 _2484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6541_ _2520_ _2524_ _2526_ _2103_ _2266_ net26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_3753_ _2853_ _2900_ _2913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4801__I B\[0\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6505__A1 _2334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6472_ _2305_ _2315_ _2455_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3684_ _1609_ _2843_ _2844_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5423_ _1282_ _1283_ _1285_ _1305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_12_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3417__I _0850_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5354_ _1228_ _1229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4305_ _0128_ _0751_ _0129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5285_ _1138_ _1150_ _1153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_99_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4236_ _3389_ _3395_ _3396_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_101_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4295__A2 _0118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4167_ _3324_ _3326_ _3327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4098_ _2958_ _2963_ _3258_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4047__A2 _3206_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6808_ _2744_ _2751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5547__A2 _1221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3558__A1 _2387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6739_ net14 _2675_ _2703_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_20_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3730__A1 _2690_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6373__I _1239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5786__A2 _1703_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3797__A1 _2886_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4210__A2 _3369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3721__A1 _2812_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5070_ _0699_ _0917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5474__A1 _3299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4021_ _3093_ _3181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5972_ _0545_ _0556_ _1907_ _1908_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4923_ _0738_ _0754_ _0755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_80_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4854_ _0617_ _0640_ _0679_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_60_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3805_ _2876_ _2890_ _2965_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4785_ _0605_ _0608_ _0609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6524_ _2500_ _2502_ _2507_ _2509_ _2510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_3736_ _2891_ _2895_ _2896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6659__S _2638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3960__A1 _3009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3667_ _2825_ _2826_ _2827_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6455_ _2044_ _2435_ _2436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5406_ _1280_ _1281_ _1284_ _1285_ _1286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6386_ _2356_ _2360_ _2361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3598_ _2277_ _2321_ _2758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_115_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3712__A1 _2858_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5337_ _0832_ _0840_ _1210_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5268_ _1131_ _1132_ _1134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4268__A2 B\[3\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5465__A1 _1293_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4219_ A\[0\]\[4\] _3379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5199_ _1057_ _1058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4706__I _0257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5768__A2 _1007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5940__A2 _0580_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6830__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5759__A2 _1596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4570_ _0314_ _2983_ _0394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3521_ _1993_ _2004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6240_ _2119_ _2200_ _2202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3452_ A\[2\]\[0\] _1246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6731__I1 _1208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6171_ _1846_ _2067_ _2126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5122_ _0886_ _0973_ _0974_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5053_ _0885_ _0896_ _0897_ _0898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5998__A2 _1208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4004_ _3161_ _3162_ _3164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4670__A2 _0492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4526__I _0282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3430__I _0850_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5955_ _0565_ _1888_ _1889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_40_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6741__I _2705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4906_ _0732_ _0735_ _0736_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5886_ _1534_ _1571_ _1814_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4837_ _0642_ _0660_ _0661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_138_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6853__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4725__A3 _0547_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4768_ _0589_ _0591_ _0592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_135_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6507_ _2361_ _2366_ _2433_ _2492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3719_ _2765_ _2879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4699_ _0345_ _0379_ _0382_ _0380_ _0523_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_140_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6438_ _2414_ _2416_ _2417_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_135_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6722__I1 _3025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6369_ _1200_ _2341_ _2342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_103_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5989__A2 _1921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5610__A1 _3351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6651__I net5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5913__A2 _0562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3924__A1 _3080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3515__I _1927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4101__A1 _3260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5601__A1 _1436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6876__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5740_ _1647_ _1652_ _1654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_43_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4955__A3 _2288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5671_ _1573_ _1577_ _1578_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4622_ _0315_ _0445_ _0446_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_129_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4553_ _0346_ _0371_ _0373_ _0375_ _0376_ _0377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_116_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3504_ _1807_ _1818_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4484_ _0307_ _2939_ _0308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5668__A1 _1504_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3435_ _1048_ _0850_ _1059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6223_ _2180_ _2182_ _2183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_143_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6154_ _2054_ _2073_ _2107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5105_ _0947_ _0950_ _0952_ _0954_ _0955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XTAP_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6085_ _1198_ _1263_ _2032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_85_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5036_ _0878_ _2922_ _2943_ _0597_ _0879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_100_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5840__A1 _1715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4643__A2 _0465_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4256__I _0079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5938_ _0303_ _0582_ _1870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6148__A2 _2046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5869_ _1762_ _1715_ _1746_ _1795_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_139_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput23 net23 result[15] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_1_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4882__A2 _0686_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6084__A1 _2027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5831__A1 _1156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4398__A1 _1301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5898__A1 _1536_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4570__A1 _0314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4322__A1 _0092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4873__A2 _0699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6841_ _0024_ net11 net1 A\[3\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_39_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6505__B _2489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4804__I _0627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4389__A1 _0200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6772_ _2645_ _3262_ _2724_ _2727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3984_ _3131_ _3142_ _3143_ _3144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5050__A2 _0608_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5723_ _1295_ _1629_ _1339_ _1635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_5654_ _1557_ _1558_ _1559_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4605_ _0419_ _0428_ _0429_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6550__A2 _2527_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5585_ _1482_ _1007_ _1309_ _1483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4561__A1 _3368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4536_ _0071_ _0353_ _3386_ _0360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_144_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6302__A2 _1811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4467_ _0202_ _0290_ _0291_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6206_ _2158_ _2163_ _2164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4313__A1 _0136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3418_ A\[3\]\[3\] _0872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4398_ _1301_ _0088_ _0222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6137_ _2049_ _2088_ _2089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5370__I _0612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6068_ _1227_ _1233_ _2013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_73_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5019_ _0790_ _0859_ _0860_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_96_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6541__A2 _2524_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4855__A2 _0629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5583__A3 _1480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6532__A2 _2513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5370_ _0612_ _1247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4321_ _0099_ _0143_ _0144_ _0145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4252_ _0075_ _1982_ _3095_ _3387_ _0076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_45_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4183_ _3339_ _3342_ _3343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__3703__I _0949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6048__A1 _1221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6599__A2 _2572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6824_ _0007_ net11 net1 A\[0\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6755_ _2671_ _2117_ _2712_ _2715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3967_ _3092_ _3125_ _3126_ _3127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4782__A1 _1356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5706_ _1352_ _1355_ _1616_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6686_ net7 _2665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3898_ _3055_ _3056_ _3058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_136_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5637_ _0230_ _0706_ _1540_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6523__A2 _2508_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5365__I _0888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4534__A1 _3096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4534__B2 _3039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5568_ _1413_ _1462_ _1463_ _1464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4519_ _2907_ _0342_ _0343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5499_ _1387_ _1388_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4837__A2 _0660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6039__A1 _1923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5262__A2 _1069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5014__A2 _0847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5317__A3 _1187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6514__A2 _2478_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4525__A1 _0331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3523__I _1147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6450__A1 _2422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5253__A2 _1112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6770__S _2724_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4870_ _0683_ _0688_ _0691_ _0695_ _0697_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_60_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5005__A2 _0803_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3821_ _2903_ _2906_ _2980_ _2981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6540_ _1786_ _1791_ _2526_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__3567__A2 _2495_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3752_ _2842_ _2846_ _2911_ _2912_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6471_ _2434_ _2436_ _2451_ _2453_ _2454_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3683_ B\[3\]\[5\] A\[3\]\[4\] _2843_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5185__I _1042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6505__A2 _2467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5422_ _1299_ _1303_ _1304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4516__A1 _0336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5353_ _0586_ _1228_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6269__A1 _2012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4304_ A\[1\]\[4\] _0128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5284_ _1137_ _1151_ _1152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4235_ _3381_ _3391_ _3394_ _3395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_68_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5492__A2 _3299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4166_ _3325_ _2310_ _3326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4097_ _3242_ _3256_ _3257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_55_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6807_ _2750_ _0059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5547__A3 _0152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4999_ _0836_ _2949_ _0837_ _1367_ _0838_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3558__A2 _2398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6738_ _2702_ _0031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6669_ _2279_ _2632_ _2650_ _0007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5180__A1 _0718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3730__A2 _2644_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5483__A2 _0770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3494__A1 _1620_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4174__I _3333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4746__A1 _0265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3518__I B\[1\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6499__A1 _2449_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3721__A2 _2806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6765__S _2719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4020_ _3167_ _3179_ _3180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_96_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5474__A2 _0600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3485__A1 _0872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4029__A3 _3186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5971_ _0551_ _0555_ _1907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_64_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4084__I _2879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4922_ _0741_ _0753_ _0754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_80_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4853_ _0642_ _0660_ _0611_ _0678_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_3804_ _2958_ _2963_ _2964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4784_ _0606_ _0595_ _0607_ _0608_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_119_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6523_ _1788_ _2508_ _2101_ _2509_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3735_ _2893_ _2894_ _2684_ _2895_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_101_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3428__I _0872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6454_ _2361_ _2366_ _2433_ _2421_ _2435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3666_ _2515_ _2484_ _2826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5405_ _0623_ _0065_ _1285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6385_ _2231_ _2358_ _2359_ _2360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3597_ _2676_ _2753_ _2757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3712__A2 _2871_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5336_ _1199_ _1208_ _1209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6675__S _2656_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5267_ _1131_ _1132_ _1133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4218_ _3329_ _3330_ _3378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_68_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5198_ _1046_ _1055_ _1056_ _1057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_29_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4149_ _3308_ _3309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6414__A1 _1975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5217__A2 _1077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4722__I _0220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4728__A1 _0133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5153__A1 _3106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4900__A1 _0626_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4900__B2 _0705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3467__A1 _1334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3801__I _1158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4719__A1 _0263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3520_ A\[2\]\[3\] _1993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3451_ _1224_ _1235_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6170_ _2112_ _2123_ _2125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_34_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5121_ _1323_ _0972_ _0973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6644__A1 _2629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5052_ _0893_ _0895_ _0897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4003_ _3161_ _3162_ _3163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_77_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5954_ _1886_ _1887_ _1888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_52_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4905_ _0733_ _0734_ _2814_ _2810_ _0735_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_80_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5885_ _1573_ _1577_ _1812_ _1813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4836_ _0648_ _0659_ _0660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_53_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5383__A1 _1219_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4767_ _0590_ _0740_ _0591_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4725__A4 _0548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6506_ _1924_ _2491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3718_ _2668_ _2876_ _2877_ _2830_ _2878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_135_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4698_ _3371_ _0242_ _0522_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5135__A1 _0983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6437_ _2415_ _2300_ _2416_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3649_ _2763_ _2809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5373__I _0733_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6368_ _2246_ _2247_ _2007_ _2341_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3697__A1 _2808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5319_ _0907_ _0942_ _1190_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6299_ _1269_ _2266_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_103_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6635__A1 _0304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5438__A2 _1319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3449__A1 _1169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5610__A2 _0951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3621__A1 _1532_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5374__A1 _1250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3924__A2 _3082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4885__B1 _0712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4101__A2 _3034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3531__I _2102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3612__A1 _1422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5670_ _1574_ _1575_ _1577_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4621_ _0432_ _0435_ _0445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4552_ _3373_ _0372_ _0371_ _0376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_117_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6510__C _1923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3503_ _1796_ _1807_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4483_ _3301_ _0307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6222_ _2181_ _2182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5668__A2 _1505_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3434_ A\[3\]\[5\] _1048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6153_ _2084_ _2085_ _2082_ _2106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6617__A1 _2147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5104_ _0953_ _2848_ _2922_ _0948_ _0954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6084_ _2027_ _2030_ _2031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5035_ _0652_ _0878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6752__I _2713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6820__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5937_ _0383_ _0514_ _0519_ _1869_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_53_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5868_ _1761_ _1781_ _1783_ _1793_ _1794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4819_ B\[2\]\[6\] _0643_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5356__A1 _2938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5799_ _0318_ _1043_ _1718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput24 net24 result[16] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_27_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6148__B _1270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6084__A2 _2030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5831__A2 _0190_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4398__A2 _0088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5595__A1 _1441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6611__B _2043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4570__A2 _2983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6843__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3833__A1 _2991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6840_ _0023_ net11 net1 A\[2\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_78_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6771_ _2726_ _0044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3983_ _3134_ _3135_ _3143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_62_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5722_ _1629_ _1630_ _1632_ _1633_ _1634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_5653_ _1441_ _1493_ _1558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4604_ _0421_ _0424_ _0427_ _0428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_5584_ _0230_ _1482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4010__A1 _3102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4535_ _0353_ _0355_ _0356_ _0358_ _0359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_116_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4561__A2 _3174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4466_ _3333_ _0773_ _0290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6205_ _2159_ _2162_ _2163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6747__I _2709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4313__A2 _1004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3417_ _0850_ _0861_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4397_ _2879_ _0220_ _0221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6136_ _2051_ _2087_ _2088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_112_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6067_ _1989_ _2011_ _2012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_86_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5018_ _0855_ _0858_ _0859_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_2506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5329__A1 _1200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6657__I _2641_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5501__A1 _1350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6866__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4855__A3 _0624_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3815__A1 _2957_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4240__A1 _3399_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4320_ _0101_ _0117_ _0144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4251_ _3393_ _0075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4182_ _3340_ _3341_ _3342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_input1_I clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4059__A1 _2904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5271__A3 _1127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6823_ _0006_ net11 net1 A\[0\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6754_ _2714_ _0037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4231__A1 _2048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3966_ _3115_ _3124_ _3126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5705_ _1353_ _1354_ _1615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6685_ _2664_ _0011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4782__A2 _0596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3897_ _3055_ _3056_ _3057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_137_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5636_ _0080_ _1278_ _1539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6678__S _2656_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4534__A2 _0354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5567_ _1394_ _1409_ _1463_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4518_ _0341_ _0342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5498_ _1369_ _1386_ _1387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_137_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4449_ _2762_ _2763_ _3390_ _0111_ _0273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_104_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6119_ _1850_ _2068_ _2069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5722__A1 _1629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6770__I0 _2642_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4289__A1 _2651_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6336__B _1900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3820_ _2912_ _2979_ _2980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4213__A1 _3322_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3751_ _2909_ _2910_ _2847_ _2911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6470_ _2145_ _2453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3682_ _2798_ _2840_ _2841_ _2842_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5421_ _1294_ _1300_ _1302_ _1303_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_64_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6761__I0 _2628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5352_ _1225_ _0859_ _1226_ _1227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4303_ _3251_ _3311_ _0127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5283_ _1138_ _1150_ _1151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4234_ _3393_ _2419_ _3394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5492__A3 _3317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4165_ A\[0\]\[1\] _3325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4096_ _3250_ _3255_ _3256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_82_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6760__I _2717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6806_ _2940_ _2640_ _2745_ _2750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4998_ _0588_ _0837_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5547__A4 _0546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5952__A1 _0075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3949_ _2931_ _3043_ _3108_ _3045_ _3109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6737_ _2673_ _2002_ _2698_ _2702_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6668_ _2649_ _2632_ _2650_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5619_ _1449_ _1461_ _1519_ _1520_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5704__A1 _1604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6599_ _1178_ _2572_ _2585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5180__A2 _0951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4691__A1 _0345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3494__A2 _0872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4443__A1 _0107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6670__I net3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6603__C _1270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4190__I A\[1\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6120__A1 _1845_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3485__A2 _1598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4365__I _3311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5970_ _1884_ _1904_ _1906_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_93_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4434__A1 _1785_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4921_ _0748_ _0752_ _0753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_64_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4852_ _0671_ _0676_ _0677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6187__A1 _2094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3803_ _2959_ _2960_ _2962_ _2963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_127_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4783_ _0600_ _0993_ _0607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6522_ _1731_ _0490_ _1772_ _0491_ _2508_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3734_ _2037_ _2894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6453_ _2421_ _2367_ _2433_ _2434_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3665_ A\[2\]\[7\] _1927_ _2825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5404_ _1282_ _1283_ _1284_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_118_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5162__A2 _1017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6384_ _2357_ _2257_ _2359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3596_ _2718_ _2746_ _2753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_127_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5335_ _3116_ _1208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3444__I B\[1\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6111__A1 _1897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5266_ _1071_ _1077_ _1063_ _1132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_4217_ _3375_ _3376_ _3377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_130_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5197_ _1047_ _1054_ _1056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5870__B1 _1794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4148_ A\[1\]\[3\] _3308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6691__S _2666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6414__A2 _1978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4079_ _3232_ _3238_ _3239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4425__A1 _0197_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4976__A2 _0766_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6178__A1 _2057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4728__A2 _2942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_78 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3951__A3 _3042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5689__B1 _3368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5153__A2 _1007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4900__A2 _0727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4113__B1 _3244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3467__A2 _1400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4664__A1 _3182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6405__A2 _2198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4185__I A\[1\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4416__A1 _0195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4967__A2 _0802_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4719__A2 _0277_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6716__I0 _2671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3450_ B\[1\]\[5\] _1224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6776__S _2724_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5120_ _0625_ _0972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5051_ _0893_ _0895_ _0896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_112_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4655__A1 _0412_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4002_ _3104_ _3112_ _3094_ _3162_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_37_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4407__A1 _0230_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5953_ _0561_ _1301_ _1887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_80_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5080__A1 _0925_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4904_ B\[0\]\[7\] _0734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5884_ _1811_ _0530_ _1578_ _1812_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_61_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5907__A1 _1562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4835_ _0654_ _0658_ _0659_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_21_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6580__A1 _0506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4766_ B\[2\]\[5\] _0590_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6505_ _2334_ _2467_ _2489_ _2490_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3717_ _2805_ _2829_ _2877_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_107_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4697_ _3371_ _0242_ _0521_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_106_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3648_ _2277_ _2805_ _2807_ _2636_ _2808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_20_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5135__A2 _0986_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6436_ _2287_ _2292_ _2415_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_136_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6367_ _2338_ _2339_ _2340_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3579_ _1993_ _1191_ _2627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3697__A2 _2816_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4894__A1 _0704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5318_ _0907_ _0942_ _1189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_88_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6298_ _2224_ _2228_ _2263_ _0585_ _2264_ _2265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_114_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6635__A2 _0525_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5249_ _1108_ _1111_ _1112_ _1113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_5_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3449__A2 _1202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6875__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5071__A1 _0917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3621__A2 _1598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6571__A1 _0506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5374__A2 _1248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4885__B2 _2452_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6866__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4620_ _0401_ _0442_ _0443_ _0444_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4551_ _0374_ _0375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3502_ _1576_ _1796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6314__A1 _2117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4482_ _3075_ _0189_ _0306_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6221_ _2148_ _2149_ _2178_ _2181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_104_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3433_ _0839_ _0894_ _0938_ _1026_ _1037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_125_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4876__A1 _0697_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6152_ _2049_ _2088_ _2105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5103_ _0946_ _0953_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6617__A2 _2602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6083_ _1204_ _2028_ _2029_ _2030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_100_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5034_ _0905_ _0829_ _0877_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6857__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5053__A1 _0885_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5936_ _3294_ _1266_ _1270_ _1868_ net19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_53_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4800__A1 _0623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5867_ _1765_ _1784_ _1792_ _1793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_139_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4818_ _0617_ _0640_ _0641_ _0642_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5356__A2 _0958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5798_ _1589_ _1716_ _1669_ _1717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_119_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4749_ _0273_ _0572_ _0573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput25 net25 result[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_6419_ _3291_ _2395_ _2396_ _2397_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_89_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6848__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5292__A1 _1154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4463__I _0286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3807__I _2190_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4858__A1 _2157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6839__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3833__A2 _2992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_0 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6770_ _2642_ _3034_ _2724_ _2726_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5586__A2 _1483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3982_ _3134_ _3135_ _3142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_51_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3597__A1 _2676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5721_ _0694_ _0220_ _0149_ _0687_ _1633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_94_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5652_ _1489_ _1492_ _1557_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4603_ _0425_ _0426_ _0427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5583_ _1478_ _1479_ _1480_ _1481_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_117_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4010__A2 _3169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4534_ _3096_ _0354_ _0357_ _3039_ _0358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_144_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4465_ _2942_ _3353_ _0289_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6204_ _3243_ _2160_ _2161_ _2162_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3416_ B\[3\]\[1\] _0850_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4396_ _3399_ _0220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5510__A2 _0594_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6135_ _2074_ _2086_ _2087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_86_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3452__I A\[2\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6066_ _1998_ _2010_ _2011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_85_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5274__A1 _3102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5017_ _0856_ _0857_ _0858_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5919_ _1549_ _1849_ _1850_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6526__A1 _1718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5329__A2 _3225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3627__I _1444_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4552__A3 _0371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4458__I _0281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3579__A1 _1993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6622__B _2597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4240__A2 _2310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6517__A1 _3103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4528__B1 _3034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3751__A1 _2909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4250_ _0073_ _2697_ _0074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4181_ A\[1\]\[3\] _1598_ _3341_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5256__A1 _1116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3806__A2 _2959_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6822_ _0005_ net11 net1 A\[0\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6753_ _2669_ _1241_ _2712_ _2714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3965_ _3115_ _3124_ _3125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4231__A2 _3390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5704_ _1604_ _1611_ _1613_ _1614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3896_ _1905_ _2576_ _3056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6684_ _2663_ _0530_ _2656_ _2664_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5635_ _1241_ _1486_ _1538_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3447__I B\[1\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5566_ _1394_ _1409_ _1462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6758__I _2716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4517_ _0318_ _0341_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5497_ _1370_ _1385_ _1386_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4448_ _2766_ _3382_ _0069_ _1290_ _0272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5495__A1 _1379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6694__S _2666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4379_ _0184_ _0202_ _0203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_98_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6118_ _1846_ _2067_ _2068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_85_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6049_ _1250_ _3263_ _1992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5798__A2 _1716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6833__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6770__I1 _3034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5722__A2 _1630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4289__A2 _0112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5486__A1 _1371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5486__B2 _1364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6617__B _2500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5410__A1 _1287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3750_ _2849_ _2910_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3972__A1 _3120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3681_ _2779_ _2795_ _2841_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5420_ _1296_ _0111_ _1302_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6761__I1 _0407_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5351_ _0855_ _0858_ _1226_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4302_ _3336_ _0098_ _0125_ _0126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5282_ _1144_ _1149_ _1150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4233_ _3392_ _3393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4164_ _3323_ _2651_ _3324_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5492__A4 _0870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4095_ _3252_ _3254_ _3255_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_95_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6805_ _2749_ _0058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4997_ _0833_ _0836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4204__A2 _3363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6856__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6736_ _2701_ _0030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3948_ _2882_ _3108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5952__A2 _2809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6667_ net10 _2649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3879_ _2113_ _3039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5618_ _1470_ _1518_ _1519_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6598_ _3206_ _2569_ _2582_ _2584_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5549_ _1439_ _1442_ _1443_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_2_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5468__A1 _0590_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4140__A1 _3299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4443__A2 _2644_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5640__A1 _1537_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3651__B1 _2810_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3954__A1 _3104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5459__A1 _1341_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5631__A1 _1496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4434__A2 _0257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4920_ _0727_ _0749_ _0750_ _0752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__6879__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4851_ _0675_ _2910_ _0676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4198__A1 _3338_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3802_ _2893_ _2961_ _2962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4782_ _1356_ _0596_ _0606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3945__A1 _2070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6521_ _0492_ _2226_ _2503_ _2506_ _1159_ _2507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_3733_ _2892_ _2893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5147__B1 _1000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6452_ _2431_ _2432_ _2433_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3664_ _2725_ _2822_ _2823_ _2824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5403_ _3399_ _0618_ _1283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3595_ _2684_ _2725_ _2739_ _2746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_6383_ _2357_ _2257_ _2358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5334_ _1205_ _1206_ _1207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6111__A2 _1229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5265_ _1129_ _1130_ _1131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4216_ _3336_ _3337_ _3376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5196_ _1047_ _1054_ _1055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_69_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4147_ _0861_ _3307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4078_ _3234_ _3237_ _3238_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_43_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6771__I _2726_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6719_ _2347_ _2679_ _2689_ _0023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5689__A1 _1595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5689__B2 _1596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4113__A1 _1312_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4664__A2 _0473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5861__A1 _1771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4416__A2 _0239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3545__I _2190_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5050_ _0605_ _0608_ _0593_ _0895_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_4001_ _3159_ _3160_ _3161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6792__S _2738_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4407__A2 _2894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5952_ _0075_ _2809_ _1886_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5080__A2 _0926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4903_ B\[0\]\[6\] _0733_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5883_ _1526_ _1811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4834_ _0650_ _0656_ _0657_ _0658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_33_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5907__A2 _1836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4765_ _1070_ _0588_ _0589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6504_ _2468_ _2466_ _2488_ _2489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3716_ _2387_ B\[1\]\[4\] _2876_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4696_ _0383_ _0514_ _0519_ _0520_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_135_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6435_ _2412_ _2413_ _2414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3647_ _2651_ _2660_ _2310_ _2806_ _2807_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6366_ _2251_ _2255_ _2339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3578_ _2376_ _2555_ _2606_ _2616_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4894__A2 _0721_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5317_ _1036_ _1183_ _1187_ _1188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__6766__I _2722_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6297_ _0685_ _2264_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5248_ _0994_ _1022_ _1112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_25_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5843__A1 _1156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5179_ _1034_ _1035_ _1036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_56_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3909__A1 _2839_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6571__A2 _2226_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4885__A2 _0686_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6087__A1 _1198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5834__A1 _1754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4270__B1 A\[0\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6360__B _2331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6562__A2 _1780_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4550_ _0340_ _0343_ _0374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4573__B2 _0384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3501_ B\[3\]\[7\] _1785_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4481_ _0971_ _3309_ _0305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6220_ _2148_ _2149_ _2178_ _2180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3432_ _0971_ _0982_ _0993_ _1015_ _1026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4876__A2 _0701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6151_ _2051_ _2087_ _2104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6078__A1 _2012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5102_ _1796_ _0951_ _0952_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6082_ _1207_ _1262_ _2029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4628__A2 _0451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5825__A1 _1715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5033_ _0651_ _0982_ _0876_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6250__A1 _2131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5935_ _1274_ _1867_ _1868_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4800__A2 _2931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5866_ _1786_ _1791_ _1792_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4817_ _0631_ _0639_ _0641_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6553__A2 _2491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5797_ _0314_ _0953_ _1716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4564__A1 _0387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4748_ _0569_ _0571_ _0572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_135_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6697__S _2666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4679_ _0469_ _0502_ _0503_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6418_ _2391_ _2394_ _2396_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_134_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput26 net26 result[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_89_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6349_ _2318_ _2217_ _2320_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4619__A2 _0441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5816__A1 _1727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5292__A2 _1142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6241__A1 _2118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6544__A2 _3191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4858__A2 _0682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3823__I _1015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5807__A1 _0980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5283__A2 _1150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4654__I _0408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3981_ _2997_ _3140_ _3141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5720_ _0065_ _0690_ _1632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5651_ _1507_ _1513_ _1555_ _1556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6535__A2 _2491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4602_ _0359_ _0360_ _0426_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5582_ _0561_ _0972_ _1480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4533_ _0149_ _0357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4464_ _0287_ _2940_ _0132_ _0288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4849__A2 _0667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6203_ _3264_ _3245_ _2161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3415_ _0817_ _0828_ _0839_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4395_ _0113_ _0217_ _0218_ _0162_ _0219_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6134_ _2084_ _2085_ _2086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_97_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6065_ _2001_ _2009_ _2010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5274__A2 _1140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5016_ _0635_ _0633_ _2267_ _2660_ _0857_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__6471__B2 _2453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6223__A1 _2180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5918_ _1221_ _0075_ _1849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4785__A1 _0605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5395__I _1273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5849_ _1772_ _3369_ _1773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4537__A1 _0359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3760__A2 _2919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5017__A2 _0857_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6214__A1 _2003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3579__A2 _1191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4528__A1 _0350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4528__B2 _0351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3751__A2 _2910_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4649__I _3369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4180_ _0773_ A\[1\]\[2\] _3340_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5256__A2 _1119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6453__A1 _2421_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6821_ _0004_ net11 net1 A\[0\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_91_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6752_ _2713_ _0036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4767__A1 _0590_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3964_ _3117_ _3120_ _3123_ _3124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__5964__B1 _1898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5703_ _1612_ _1156_ _1607_ _1610_ _1613_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6683_ net6 _2663_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3895_ _3031_ _3053_ _3054_ _3055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4519__A1 _2907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5634_ _1423_ _1424_ _1481_ _1483_ _1537_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3990__A2 _3145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5192__A1 _3081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5192__B2 _1042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5565_ _1459_ _1460_ _1461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_129_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4516_ _0336_ _0339_ _0340_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5496_ _1374_ _1377_ _1384_ _1385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_144_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4447_ _0160_ _0265_ _0270_ _0232_ _0271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3463__I _1356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4378_ A\[1\]\[5\] B\[3\]\[4\] _0202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6117_ _1849_ _2066_ _2067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6048_ _1221_ _3269_ _1991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4930__A1 _0730_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5486__A2 _1372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5410__A2 _1288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3548__I B\[1\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3680_ _2779_ _2795_ _2840_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_118_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5350_ _0824_ _1223_ _3246_ _3247_ _1225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_86_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4301_ _0091_ _0097_ _0125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5281_ _1146_ _1148_ _1149_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5477__A2 _0599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4232_ A\[0\]\[5\] _3392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4163_ A\[0\]\[2\] _3323_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5229__A2 _1089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4094_ _2946_ _3253_ _3254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_83_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6543__B _2226_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3660__A1 _2676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6804_ _3174_ _2637_ _2745_ _2749_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4996_ _0766_ _0834_ _0835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5401__A2 _0620_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6735_ _2671_ _2003_ _2698_ _2701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3947_ _3039_ _3106_ _3107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3412__A1 _0729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3458__I _1301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6666_ _2648_ _0006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3878_ _3037_ _2806_ _3038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5165__A1 _0913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6769__I _2717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5617_ _1472_ _1517_ _1518_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6597_ _3206_ _2569_ _2582_ _2583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5548_ _1434_ _1440_ _1441_ _1442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5479_ _1362_ _1365_ _1366_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__3479__A1 _1081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4140__A2 _0751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3921__I _1576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6417__A1 _2391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output26_I net26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3651__A1 _2809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5848__I _0980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6453__B _2433_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3651__B2 _1301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3954__A2 _3112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5156__A1 _1003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3890__A1 _3047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4850_ B\[2\]\[7\] _0675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3801_ _1158_ _2961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4198__A2 _3356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4781_ _0595_ _0598_ _0601_ _0604_ _0605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_6520_ _2368_ _2504_ _2506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3732_ A\[2\]\[7\] _2892_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3945__A2 _2026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5147__A1 _2933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6451_ _2422_ _2423_ _2429_ _2432_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_119_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3663_ _2732_ _2821_ _2168_ _2398_ _2823_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_9_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5147__B2 _3035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5402_ _0161_ _0625_ _1282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6382_ _2235_ _2357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3594_ _2732_ _2168_ _2739_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5333_ _0819_ _0865_ _1206_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5264_ _1062_ _2849_ _1130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6538__B _1273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4215_ _3327_ _3331_ _3375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5195_ _1052_ _1053_ _1054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_69_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4146_ _2863_ _3305_ _3306_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3881__A1 _3039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6823__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4077_ _2929_ _3235_ _3236_ _3237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5386__A1 _1198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4979_ _0812_ _0815_ _0816_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_138_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6718_ _2649_ _2679_ _2689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6649_ _0350_ _2634_ _2632_ _2635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5689__A2 _0318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6638__A1 _2623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5310__A1 _1119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5377__A1 _0798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5377__B2 _0849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5129__A1 _0979_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5301__A1 _1123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6846__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4000_ _3093_ _2849_ _3160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5604__A2 _3313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5951_ _0566_ _0573_ _1885_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4812__B1 _2814_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4902_ _0731_ _2354_ _2026_ _0612_ _0732_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5882_ _1528_ _1582_ _1810_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5368__A1 _0847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4833_ _2787_ _0599_ _0657_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4764_ B\[2\]\[4\] _0588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6503_ _2308_ _2486_ _2465_ _2487_ _2488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3715_ _2818_ _2833_ _2874_ _2875_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4695_ _0515_ _0518_ _0519_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_101_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6434_ _2407_ _2410_ _2405_ _2413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3646_ _2190_ _2806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5540__A1 _1248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6365_ _2237_ _2250_ _2338_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3577_ _2473_ _2545_ _2606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5316_ _1184_ _1186_ _1187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_115_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6296_ _2230_ _2262_ _2263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_130_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5247_ _1097_ _1109_ _1110_ _1111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_64_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5843__A2 _0190_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5178_ _0940_ _0941_ _0907_ _1035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_111_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6782__I _2734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4129_ net15 _3289_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5359__A1 _1227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3909__A2 _2902_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4031__A1 _3189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3646__I _2190_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5531__A1 _0079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6869__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6087__A2 _1263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4098__A1 _2958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5101__I _0600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4270__A1 _2763_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4270__B2 _2762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5770__A1 _1682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4573__A2 _0394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3500_ _1752_ _1763_ _1774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4480_ _0303_ _0304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_128_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3431_ _1004_ _1015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5522__A1 _1394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6150_ _2101_ _2103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5101_ _0600_ _0951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6081_ _1207_ _1262_ _2028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4089__A1 _2966_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5032_ _0869_ _0874_ _0875_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_111_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3836__A1 _2994_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5589__A1 _1486_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5589__B2 _0999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6250__A2 _2172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5934_ _1806_ _1866_ _1867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_40_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5865_ _1718_ _1789_ _1790_ _1791_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4850__I B\[2\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4816_ _0631_ _0639_ _0640_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_22_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5796_ _1702_ _1703_ _1678_ _1715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_119_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4747_ _0233_ _0560_ _0570_ _0266_ _0571_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4564__A2 _3075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4678_ _0480_ _0485_ _0471_ _0502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6417_ _2391_ _2394_ _2395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3629_ _2784_ _1059_ _1543_ _2788_ _2789_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__5513__A1 _0136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput27 net27 result[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_1_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6348_ _2318_ _2217_ _2319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6279_ _2238_ _2243_ _2244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_130_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3827__A1 _1796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6241__A2 _2198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4252__A1 _0075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4252__B2 _3387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5752__A1 _3367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5807__A2 _0257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3818__A1 _2925_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4491__A1 _2948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3980_ _3129_ _3130_ _3140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4243__A1 _3382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5991__A1 _0696_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5650_ _1509_ _1512_ _1555_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4601_ _0330_ _0352_ _0425_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5581_ _0623_ _0070_ _1479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4546__A2 _0368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4532_ _0281_ _3098_ _0356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4463_ _0286_ _0287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6202_ _3270_ _2160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3414_ A\[3\]\[4\] _0828_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4394_ _0148_ _0160_ _0218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_125_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6133_ _0669_ _1612_ _2085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6064_ _2006_ _2008_ _2009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5015_ _0734_ _2967_ _2092_ _0733_ _0856_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4845__I _0668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4482__A1 _3075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6223__A2 _2182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4234__A1 _3393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5917_ _1247_ _1486_ _1437_ _1222_ _1848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4785__A2 _0608_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5848_ _0980_ _1772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6526__A3 _1788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4537__A2 _0360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5779_ _1691_ _1694_ _1696_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6462__A2 _2385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6214__A2 _2172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5973__A1 _0290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4490__I _0307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5725__A1 _1634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4528__A2 _3032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4700__B3 _0518_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5256__A3 _1120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4464__A1 _0287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6820_ _0003_ net11 net1 A\[0\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_90_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6751_ _2665_ _1000_ _2712_ _2713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3963_ _3121_ _3122_ _3123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5964__A1 _1897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4767__A2 _0740_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5964__B2 _1564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5702_ _0326_ _1612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6682_ _2662_ _0010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3894_ _3051_ _3052_ _3054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5633_ _1485_ _1494_ _1535_ _1536_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5716__A1 _1607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4519__A2 _0342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5564_ _1392_ _1448_ _1460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_117_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5192__A2 _0878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4515_ _0337_ _0338_ _0339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5495_ _1379_ _1383_ _1384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4446_ _0217_ _0233_ _0270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_105_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4377_ _1565_ _3308_ _0201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6116_ _1250_ _0562_ _2066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6047_ _1245_ _1256_ _1990_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5955__A1 _0565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3919__I _2996_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6755__I0 _2671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4930__A2 _0736_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4446__A1 _0217_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5946__A1 _0537_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3829__I _1015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6746__I0 _2661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6371__A1 _2342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4921__A2 _0752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4300_ _3343_ _0122_ _0123_ _0124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5280_ _1139_ _1143_ _1148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4231_ _2048_ _3390_ _3391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4162_ _3304_ _3320_ _3321_ _3322_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4093_ _2937_ _2950_ _3253_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6803_ _2748_ _0057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4995_ _0833_ _2785_ _0834_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6734_ _2700_ _0029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3946_ _2354_ _3106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3877_ _2398_ _3037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6665_ _2119_ _2647_ _2631_ _2648_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6737__I0 _2673_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5616_ _1496_ _1516_ _1517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6362__A1 _2323_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6596_ _3147_ _3209_ _2582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4912__A2 _2821_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5547_ _1250_ _1221_ _0152_ _0546_ _1441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_133_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6114__A1 _2057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5478_ _1363_ _1358_ _1364_ _1365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_132_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4429_ _0251_ _0252_ _0253_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3479__A2 _1532_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6417__A2 _2394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4979__A2 _0815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3651__A2 _2354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output19_I net19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3649__I _2763_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6728__I0 _2663_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3890__A2 _3048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5919__A1 _1549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3559__I _2102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3800_ _1224_ _2704_ _2960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4780_ _0602_ _0603_ _0604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_53_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3731_ _2876_ _2889_ _2890_ _2891_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__6820__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3662_ _2732_ _2168_ _1938_ _2821_ _2822_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5147__A2 _0998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6450_ _2422_ _2423_ _2429_ _2431_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5401_ A\[0\]\[2\] _0620_ _1281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6381_ _2337_ _2355_ _2356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_3593_ A\[2\]\[7\] _2732_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5332_ _0821_ _0864_ _1205_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5263_ _1067_ _1128_ _1129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_138_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4658__A1 _0394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4214_ _3373_ _3374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5194_ _0876_ _1049_ _0952_ _1053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_4145_ A\[1\]\[4\] _3305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4076_ _2936_ _2954_ _3236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_83_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5083__A1 _0704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5386__A2 _1263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4978_ _0813_ _0814_ _0815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6717_ _2688_ _0022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3929_ _3078_ _3087_ _3088_ _3089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_50_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6648_ net4 _2634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6579_ _0506_ _0507_ _0510_ _2564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_124_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4897__A1 _0634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_35 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5310__A2 _1120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6878__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5074__A1 _0915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3624__A2 _0949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4821__A1 _0588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5377__A2 _1240_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5129__A2 _0980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6869__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5950_ _0557_ _0575_ _1882_ _1884_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4812__A1 _0633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4812__B2 _0635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4901_ _0633_ _0731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5881_ _1529_ _1808_ _1581_ _1809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4832_ _2790_ _0655_ _0656_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6565__A1 _1793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5368__A2 _1243_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4763_ _0586_ _1796_ _0587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6502_ _2458_ _2461_ _2487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3714_ _2820_ _2832_ _2874_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4694_ _0454_ _0516_ _0517_ _0518_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6433_ _2406_ _2411_ _2412_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3645_ _2495_ _2299_ _2805_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3576_ _1905_ _2576_ _2586_ _2596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6364_ _2252_ _2254_ _2337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6549__B _2533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5540__A2 _0281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5315_ _1116_ _1181_ _1185_ _1186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6295_ _2258_ _2261_ _2262_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5246_ _1100_ _1101_ _1110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_102_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5177_ _0991_ _1032_ _1033_ _1034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4128_ net16 _3288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4583__I _3101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4059_ _2904_ _2905_ _2903_ _3219_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6556__A1 _1981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3909__A3 _2904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6308__A1 _1526_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5531__A2 _1296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3542__A1 _2135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4098__A2 _2963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5047__A1 _0889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4493__I _2948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4270__A2 A\[0\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6213__I _2907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5770__A2 _1683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3781__A1 _2938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3430_ _0850_ _1004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3533__A1 _1960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5100_ _0948_ _2848_ _0950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6080_ _1985_ _2025_ _2027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5286__A1 _1073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5031_ _0871_ _0873_ _0874_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3836__A2 _2995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5589__A2 _0998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5933_ _1864_ _1865_ _1866_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4261__A2 _0084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6538__A1 _3191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5864_ _1787_ _1788_ _1790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4815_ _0637_ _0638_ _0639_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5210__A1 _1065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5795_ _1662_ _1713_ _1714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4013__A2 _3172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4746_ _0265_ _0267_ _0570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_119_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5962__I _0287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4677_ _0460_ _0468_ _0501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6416_ _1935_ _1979_ _2183_ _2393_ _2182_ _2394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__5513__A2 _0655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3628_ _2785_ _0861_ _2786_ _2787_ _2788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput17 net17 result[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput28 net28 result[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_6347_ _2194_ _2318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3559_ _2102_ _2419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6278_ _2239_ _2242_ _2243_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5229_ _1080_ _1089_ _1091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3827__A2 _0927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5029__A1 _2984_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5202__I _0969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4252__A2 _1982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6529__A1 _1044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6836__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5752__A2 _1043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6701__A1 _2629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4491__A2 _0313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5112__I _0836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4243__A2 _1158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5440__A1 _1307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4600_ _0329_ _0422_ _0423_ _0424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5580_ _1311_ _1278_ _1478_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4531_ _3101_ _0354_ _0355_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4462_ A\[1\]\[7\] _0286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6201_ _1239_ _3243_ _2159_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3506__A1 _1785_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3413_ B\[3\]\[2\] _0817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4393_ _0072_ B\[1\]\[4\] _0217_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6132_ _2082_ _2083_ _2084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6063_ _0834_ _2007_ _2008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5014_ _0749_ _0847_ _0854_ _0797_ _0855_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_38_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4482__A2 _0189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6759__A1 _2654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4234__A2 _2419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4861__I _0686_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6859__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5916_ _1843_ _1844_ _1846_ _1847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_35_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3993__A1 _3148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5847_ _1732_ _1770_ _1771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5778_ _1691_ _1694_ _1695_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3745__A1 _2839_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4729_ _0286_ _0751_ _0553_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5498__A1 _1369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4170__A1 _3324_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5422__A1 _1299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5725__A2 _1635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5489__A1 _1375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4464__A2 _2940_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6750_ _2705_ _2712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_51_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3962_ _3047_ _3048_ _3122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5964__A2 _0317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3975__A1 _3031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5701_ _1608_ _1610_ _1611_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_31_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6681_ _2661_ _0191_ _2656_ _2662_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3893_ _3051_ _3052_ _3053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5632_ _1476_ _1484_ _1535_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5563_ _1457_ _1458_ _1459_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4514_ _3298_ _3303_ _0338_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5494_ _1381_ _1382_ _1383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_117_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4445_ _0264_ _0268_ _0269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_144_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4152__A1 _3311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4376_ _0147_ _0198_ _0199_ _0200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6115_ _1847_ _1855_ _2065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6046_ _1236_ _1259_ _1988_ _1989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5404__A1 _1282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5687__I _0963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6601__B1 _2587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3966__A1 _3115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6879_ _0062_ net11 net1 B\[3\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_10_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6755__I1 _2117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3935__I _3037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6380__A2 _2353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5643__A1 _0561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4446__A2 _0233_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5643__B2 _1311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6691__I0 _2669_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3957__A1 _3006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6746__I1 _1007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3845__I _3004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4382__A1 _0136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4134__A1 _0696_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4230_ A\[0\]\[3\] _3390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5882__A1 _1528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4161_ _3315_ _3319_ _3321_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4092_ _3251_ _2949_ _3252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5634__A1 _1423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5634__B2 _1483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6802_ _3075_ _2634_ _2745_ _2748_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5937__A2 _0514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4994_ B\[2\]\[5\] _0833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6733_ _2669_ _0979_ _2698_ _2700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3945_ _2070_ _2026_ _3105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6664_ net9 _2647_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3876_ _2932_ _3032_ _3034_ _3035_ _3036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6737__I1 _2002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5615_ _1498_ _1515_ _1516_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_104_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6595_ _0452_ _0459_ _2580_ _2581_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_118_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5546_ _1247_ _0546_ _1440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4912__A3 _0716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5477_ A\[1\]\[3\] _0599_ _1364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4428_ _0201_ _0203_ _0252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4359_ _0124_ _0181_ _0182_ _0183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5625__A1 _1526_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6029_ _0979_ _2908_ _1970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6728__I1 _3225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6353__A2 _0524_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4364__A1 _0183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5616__A1 _1496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5120__I _0625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5919__A2 _1849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6041__A1 _1526_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3730_ _2690_ _2644_ _2890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5276__B _1142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3661_ A\[2\]\[6\] _2821_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5400_ _0149_ _1278_ _1280_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6380_ _2340_ _2353_ _2355_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3592_ _2146_ _2484_ _2725_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5331_ _1203_ _1204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4107__A1 _2959_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5262_ _1065_ _1069_ _1128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_142_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4213_ _3322_ _3357_ _3373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5193_ _1049_ _1050_ _1051_ _1038_ _1052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_69_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4144_ _3298_ _3303_ _3304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_56_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5607__A1 _1503_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4075_ _2936_ _2954_ _3235_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_55_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5083__A2 _0721_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6280__A1 _1244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4977_ _0765_ _0767_ _0814_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6716_ _2671_ _2240_ _2678_ _2688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3928_ _3079_ _3086_ _3088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6647_ _2633_ _0000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3859_ _0729_ _0795_ _3019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4346__A1 _0107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6578_ _1794_ _1795_ _2563_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_118_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5529_ _1419_ _1316_ _1420_ _1421_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6099__A1 _1811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5846__A1 _1683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6646__I0 _0490_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5074__A2 _0918_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4821__A2 _1532_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6023__A1 _3250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4585__A1 _0406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3609__B _2761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5129__A3 _0975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6262__A1 _3295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4812__A2 _1246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4900_ _0626_ _0727_ _0728_ _0705_ _0730_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_46_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5880_ _1470_ _1518_ _1808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_61_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4831_ B\[2\]\[1\] _0655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6565__A2 _1781_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4762_ B\[2\]\[6\] _0586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4040__A3 _3194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6501_ _2458_ _2461_ _2486_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3713_ _2855_ _2872_ _2873_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4693_ _0457_ _0458_ _0517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6432_ _2407_ _2410_ _2411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3644_ _2764_ _2803_ _2804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6363_ _1925_ _2334_ _2335_ _2336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3575_ _2256_ _2565_ _2586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5314_ _1119_ _1120_ _1185_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_114_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6294_ _2259_ _2260_ _2261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5828__A1 _1717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5245_ _1100_ _1101_ _1109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_130_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5176_ _1030_ _1031_ _1033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6565__B _0696_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4864__I _0689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4127_ _3224_ _3286_ _3287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4058_ _2906_ _3068_ _3216_ _3217_ _3211_ _3213_ _3218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai33_1
XFILLER_24_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6800__I0 _0472_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4567__A1 _0387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6308__A2 _2273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4319__A1 _0101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4104__I _3263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3542__A2 _2223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6492__A1 _2275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6244__A1 _0565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6547__A2 _2368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4014__I _3072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5507__B1 _3313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3781__A2 _2940_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4730__A1 _0290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5286__A2 _1141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5030_ _0833_ _1576_ _0873_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4797__A1 _2882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5932_ _1809_ _1810_ _1863_ _1865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_81_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5863_ _1787_ _1788_ _1789_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4814_ _0634_ _0636_ _0632_ _0638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5794_ _1663_ _1706_ _1709_ _1711_ _1712_ _1713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_21_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5210__A2 _1067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4745_ _0567_ _0568_ _0569_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4676_ _0401_ _0431_ _0441_ _0500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__4859__I B\[0\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6415_ _2392_ _2180_ _2393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3627_ _1444_ _2787_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3763__I _2922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput18 net18 result[10] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_66_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput29 net29 result[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_6346_ _2302_ _2316_ _2317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_3558_ _2387_ _2398_ _2408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6277_ _2115_ _2160_ _2241_ _2242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3489_ _1587_ _1642_ _1653_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_88_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5228_ _1080_ _1089_ _1090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4485__B1 _0256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5159_ _1011_ _1012_ _1014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5029__A2 _0870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3460__A1 _1312_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3938__I _2048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_122_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6217__A1 _2173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4491__A3 _0314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4228__B1 _3387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4009__I _3096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4779__A1 _0594_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5440__A2 _1322_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3848__I _1246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4530_ _3385_ _0354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4951__A1 _0727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4461_ _0283_ _0221_ _0225_ _0284_ _0285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_116_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3583__I _1949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6200_ _3266_ _1948_ _2158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4703__A1 _0304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3506__A2 _1829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3412_ _0729_ _0795_ _0806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4392_ _0157_ _0174_ _0215_ _0216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5900__B1 _1560_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6131_ _2077_ _2080_ _2083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5259__A2 _1089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6062_ _2005_ _1955_ _2007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5013_ _0785_ _0798_ _0854_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_39_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6208__A1 _3275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3690__A1 _1785_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5431__A2 _1309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5915_ _1539_ _1845_ _1846_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5846_ _1683_ _1769_ _1770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5195__A1 _1052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5777_ _1692_ _1693_ _1694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4728_ _0133_ _2942_ _0552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4942__A1 _1499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3745__A2 _2902_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4659_ _3182_ _3369_ _0479_ _0483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_66_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6329_ _2293_ _2295_ _2297_ _2298_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__4170__A2 _3326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3681__A1 _2779_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5422__A2 _1303_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5369__B _1244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3433__B2 _1026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5186__A1 _2998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5883__I _1526_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4933__A1 _1444_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3617__B _2776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5489__A2 _1371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6438__A1 _2414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5110__A1 _2994_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5661__A2 _1566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6610__A1 _1183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5413__A2 _0681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3961_ _3010_ _3036_ _3121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3424__A1 _0905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5700_ _1357_ _1366_ _1610_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_17_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6680_ net5 _2661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3892_ _1916_ _2234_ _3052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5631_ _1496_ _1516_ _1533_ _1534_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5177__A1 _0991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3727__A2 _2827_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4924__A1 _0724_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5562_ _0668_ _0473_ _1458_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4513_ _3300_ _3302_ _0337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5493_ _1380_ _0392_ _0255_ _0837_ _1382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_105_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4444_ _0265_ _0266_ _0267_ _0268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_144_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4152__A2 _0927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4375_ _0151_ _0155_ _0199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6429__A1 _2272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6114_ _2057_ _2063_ _2064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_98_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6045_ _1238_ _1258_ _1988_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6826__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5652__A2 _1492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6573__B _2418_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6601__A1 _1981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5404__A2 _1283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6601__B2 _2225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3415__A1 _0817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3966__A2 _3124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6878_ _0061_ net11 net1 B\[3\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_22_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6799__I _2744_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5829_ _1722_ _1750_ _1751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4391__A2 _0173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5208__I _0917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4112__I _3271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6668__A1 _2649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5340__A1 _0827_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6691__I1 _1612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3957__A2 _3116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4382__A2 _3333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5118__I _0615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4022__I _3181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3590__B1 _2697_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4134__A2 _3293_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6849__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4160_ _3315_ _3319_ _3320_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_122_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3893__A1 _3051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4091_ _0707_ _3251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5634__A2 _1424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3645__A1 _2495_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6393__B _2368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6824__D _0007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6801_ _2747_ _0056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4993_ _0643_ _2943_ _0832_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6732_ _2699_ _0028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3944_ _3097_ _3100_ _3103_ _3104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__4070__A1 _2925_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6663_ _2646_ _0005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3875_ _1323_ _3035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5614_ _1502_ _1514_ _1515_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6594_ _2579_ _2566_ _2580_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5545_ _1282_ _1427_ _1438_ _1319_ _1439_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_117_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5028__I B\[2\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4912__A4 _0682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5476_ A\[1\]\[5\] _0655_ _1363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4867__I _0692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4427_ _0184_ _0202_ _0251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5322__A1 _0868_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3771__I _2814_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5873__A2 _1798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4676__A3 _0441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4358_ _0126_ _0141_ _0182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_59_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4289_ _2651_ _0112_ _0113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5625__A2 _0191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6028_ _1965_ _1968_ _1969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__3636__A1 _1488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3939__A2 _3098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3946__I _2354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4364__A2 _0187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4116__A2 _3275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5313__A1 _0991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5864__A2 _1788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6041__A2 _1208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3660_ _2676_ _2753_ _2819_ _2820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4355__A2 _0177_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3591_ _2179_ _2684_ _2711_ _2505_ _2718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_127_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3563__B1 _2070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5330_ _0812_ _0815_ _1201_ _1203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5261_ _1041_ _1126_ _1127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_48_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4212_ _3366_ _3370_ _3372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_142_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5192_ _3081_ _0878_ _2848_ _1042_ _1051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3866__A1 _2921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4143_ _3300_ _3302_ _3303_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_68_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4074_ _2947_ _3233_ _3234_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3618__A1 _2759_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4291__A1 _1235_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4976_ _0664_ _0766_ _0813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6715_ _2687_ _0021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4371__B _0194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4594__A2 _0416_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3927_ _3079_ _3086_ _3087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6646_ _0490_ _2628_ _2632_ _2633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3858_ _0762_ _0784_ _3018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4346__A2 _0079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6577_ _2554_ _2560_ _2562_ net29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3789_ _2787_ _2949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5528_ _0229_ _0168_ _1310_ _1002_ _1420_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_30_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6099__A2 _1817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5459_ _1341_ _1342_ _1344_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6646__I1 _2628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3609__A1 _2764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4282__A1 _0072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output24_I net24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4585__A2 _0408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5534__A1 _0112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6262__A2 _2225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4830_ _0650_ _0602_ _0607_ _0653_ _0654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XTAP_2480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4025__A1 _3024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6565__A3 _2550_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4761_ _0584_ _0585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3712_ _2858_ _2871_ _2872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6500_ _2395_ _2448_ _2483_ _2485_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4692_ _0457_ _0458_ _0516_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3643_ _2761_ _2764_ _2767_ _2803_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5525__A1 _1314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6431_ _2409_ _2286_ _2410_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6362_ _2323_ _2333_ _2335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3574_ _2256_ _2565_ _2576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_115_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5313_ _0991_ _1032_ _1184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6293_ _1985_ _2025_ _2260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5828__A2 _1720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5244_ _0962_ _1107_ _1108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3839__A1 _2948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3839__B2 _2995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5175_ _1030_ _1031_ _1032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_57_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4126_ _3228_ _3231_ _3285_ _3286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_83_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4057_ _3027_ _3066_ _3069_ _3067_ _3217_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_37_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6005__A2 _3244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4016__A1 _3082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6800__I1 _2628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4567__A2 _0319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4959_ _0744_ _0747_ _0794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4319__A2 _0117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6629_ _2603_ _2612_ _2615_ net33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5507__A1 _0836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5507__B2 _0837_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5931_ _1809_ _1810_ _1863_ _1864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4797__A2 _0620_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5994__A1 _3224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5862_ _1731_ _0476_ _1772_ _0342_ _1788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4813_ _0632_ _0634_ _0636_ _0637_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__6794__I0 _2005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5793_ _1600_ _1602_ _1676_ _1712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5210__A3 _1069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4744_ _0073_ _2969_ _2766_ _3380_ _0568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_108_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4675_ _0470_ _0498_ _0499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_119_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3626_ _0817_ _2786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6414_ _1975_ _1978_ _2392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_116_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput19 net19 result[11] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_3557_ B\[1\]\[1\] _2398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6345_ _2305_ _2315_ _2316_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_115_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6276_ _1223_ _2240_ _2241_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3488_ _1609_ _1631_ _1642_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_115_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5227_ _1082_ _1085_ _1088_ _1089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_131_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4485__A1 _0189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4485__B2 _2983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5682__B1 _0256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5158_ _1011_ _1012_ _1013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4109_ _2704_ _3269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4237__A1 _3389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5089_ _0935_ _0936_ _0937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_44_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5985__A1 _1876_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6785__I0 _1039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4960__A2 _0752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4491__A4 _2995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4228__B2 _1982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4779__A2 _0828_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6776__I0 _2673_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3864__I _2998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4460_ _0219_ _0224_ _0284_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3411_ _0762_ _0784_ _0795_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_132_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4703__A2 _0525_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4391_ _0159_ _0173_ _0215_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6130_ _2077_ _2080_ _2082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_112_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6061_ _1595_ _2002_ _2003_ _2005_ _2006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5012_ _0846_ _0852_ _0853_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_79_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3690__A2 _2849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5914_ _0888_ _1482_ _1845_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5719__A1 _0917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6767__I0 _2640_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5845_ _0476_ _1140_ _1769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3993__A3 _3152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5195__A2 _1053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5776_ _1634_ _1635_ _1693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4727_ _0549_ _0275_ _0550_ _0551_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4942__A2 B\[2\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6150__I _2101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4658_ _0394_ _0481_ _0461_ _0482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3609_ _2764_ _2767_ _2761_ _2769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4589_ _0411_ _3043_ _0354_ _3039_ _0413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6328_ _2140_ _2296_ _2297_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6259_ _2218_ _2221_ _2222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_88_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5186__A2 _1043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4933__A2 B\[2\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6060__I _1229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4697__A1 _3371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6438__A2 _2416_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4449__A1 _2762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5110__A2 _0959_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3672__A2 _2831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5949__A1 _0559_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6610__A2 _1187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3960_ _3009_ _3118_ _3119_ _3120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3424__A2 _0927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3891_ _3011_ _3036_ _3049_ _3050_ _3051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__6850__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5630_ _1473_ _1531_ _1495_ _1533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4924__A2 _0755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5561_ _1454_ _1456_ _1457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6126__A1 _1830_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4512_ _0324_ _0334_ _0335_ _0336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5492_ _1380_ _3299_ _3317_ _0870_ _1381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_144_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4443_ _0107_ _2644_ _0267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4374_ _0151_ _0155_ _0198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6113_ _2060_ _2062_ _2063_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6429__A2 _2285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6044_ _1217_ _1261_ _1986_ _1987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3663__A2 _2821_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6601__A2 _2583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3415__A2 _0828_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6877_ _0060_ net11 net1 B\[3\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__6841__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5168__A2 _1022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5828_ _1717_ _1720_ _1750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4915__A2 _0689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5759_ _0387_ _1596_ _1673_ _1674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_124_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6117__A1 _1849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6668__A2 _2632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5340__A2 _0842_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4851__A1 _0675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6832__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6356__A1 _1921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5159__A2 _1012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4382__A3 _1004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3590__A1 _2690_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3590__B2 _2704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3893__A2 _3052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4090_ _3248_ _2972_ _3249_ _3250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5095__A1 _0907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3645__A2 _2299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3589__I _2146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6800_ _0472_ _2628_ _2745_ _2747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5398__A2 _1276_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4992_ _2938_ _0830_ _0650_ _0831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_56_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6731_ _2665_ _1208_ _2698_ _2699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3943_ _3101_ _3102_ _3103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6823__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6840__D _0023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6662_ _2118_ _2645_ _2638_ _2646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3874_ _3033_ _3034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5613_ _1507_ _1513_ _1514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6593_ _0508_ _0509_ _2579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5544_ _0972_ _1437_ _0999_ _0357_ _1438_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_129_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5475_ _1358_ _1359_ _1360_ _1361_ _1362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_144_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4426_ _0200_ _0212_ _0249_ _0250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5044__I _0848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4357_ _0126_ _0141_ _0181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_28_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4288_ _0111_ _0112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6027_ _1966_ _1967_ _1968_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3636__A2 _1554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4061__A2 _3218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6338__A1 _2172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5010__A1 _2893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3572__A1 _2473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6510__A1 _2424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5077__A1 _0921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5889__I _0420_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6714__S _2682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6577__A1 _2554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4742__B _0565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4052__A2 _3152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3590_ _2690_ _2102_ _2697_ _2704_ _2711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5552__A2 _1446_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3563__A1 _2452_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3563__B2 _2430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3872__I _2961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5304__A2 _1113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5260_ _1045_ _1126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4211_ _3366_ _3370_ _3364_ _3371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_130_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5191_ _1042_ _3081_ _1050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3866__A2 _3025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4142_ _2945_ _3301_ _3302_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5068__A1 _0889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3821__B _2980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4073_ _2944_ _2952_ _3233_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4291__A2 _0114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4208__I _3367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4975_ _0764_ _0779_ _0811_ _0812_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4043__A2 _3194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6714_ _2669_ _2160_ _2682_ _2687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3926_ _3084_ _3085_ _3086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_137_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6645_ _2631_ _2632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3857_ _3003_ _3014_ _3016_ _3017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6576_ _1274_ _2561_ _2546_ _2562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4346__A3 _2102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6740__A1 _2629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3788_ _0773_ _2948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3554__A1 _2343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5527_ _0229_ _1310_ _0712_ _0168_ _1419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3782__I _1565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6298__C _2264_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5458_ _1341_ _1342_ _1343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_133_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4409_ _0102_ B\[1\]\[3\] _0233_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5389_ net2 _1267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3609__A2 _2767_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4806__A1 _0626_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4282__A2 _2484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output17_I net17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5231__A1 _1052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6839__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5782__A2 _1699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5534__A2 _0628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6798__A1 _1267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4025__A2 _3181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4760_ _3295_ _0674_ _0584_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3711_ _2862_ _2870_ _2871_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3784__A1 _2942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4691_ _0345_ _0379_ _0515_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_105_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6430_ _2269_ _2409_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3642_ _2772_ _2800_ _2801_ _2802_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5525__A2 _1317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6399__B _1957_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6361_ _2323_ _2333_ _2334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3573_ _2376_ _2555_ _2565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5312_ _1122_ _1177_ _1179_ _1182_ _1183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_6292_ _1987_ _2024_ _2259_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5289__A1 _1156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5243_ _1095_ _1096_ _1107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3839__A2 _2998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5174_ _0908_ _0937_ _1031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_111_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4125_ _3239_ _3284_ _3285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_57_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4056_ _2904_ _2905_ _3216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3777__I _2790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5213__A1 _1009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4958_ _0735_ _0792_ _0793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_51_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3909_ _2839_ _2902_ _2904_ _3069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_138_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4889_ _2892_ _0716_ _0717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6628_ _1274_ _2614_ _2546_ _2615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6559_ _3193_ _2541_ _2543_ _2500_ _2544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_106_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5452__A1 _0692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4558__A3 _3371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5755__A2 _1667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5507__A2 _3309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5443__A1 _1281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6640__B1 _2620_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5930_ _1813_ _1861_ _1863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_65_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5994__A2 _3286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5861_ _1771_ _1773_ _1787_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_61_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4812_ _0633_ _1246_ _2814_ _0635_ _0636_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_34_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5792_ _1706_ _1710_ _1711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6794__I1 _2647_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3757__A1 _2843_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4743_ _3393_ _2812_ _2813_ _0112_ _0567_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4674_ _0487_ _0497_ _0498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6413_ _2386_ _2390_ _2391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_134_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3625_ _1499_ _2785_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6344_ _2309_ _2314_ _2315_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3556_ A\[2\]\[5\] _2387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6275_ _3264_ _2240_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3487_ _1620_ _0740_ _1631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5226_ _1086_ _1087_ _1088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5682__A1 _0395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4485__A2 _3072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5682__B2 _1042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5157_ _0688_ _1003_ _0919_ _1012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_99_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4108_ _3261_ _3265_ _3267_ _3268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5088_ _0678_ _0756_ _0936_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input16_I sel_out[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5434__A1 _1309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4237__A2 _3395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4039_ _3193_ _3198_ _3199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_71_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5985__A2 _1921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6785__I1 _2637_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5936__B _1270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6162__A2 _2115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4131__I _3290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3920__A1 _2984_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4476__A2 _0299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6058__I _1955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3987__A1 _3139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6722__S _2692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5728__A2 _1639_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6776__I1 _2200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4164__A1 _3323_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3410_ _0773_ A\[3\]\[1\] _0784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4390_ _0197_ _0213_ _0214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5900__A2 _1511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3911__A1 _0718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3880__I _2810_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6060_ _1229_ _2005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input8_I input_val[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5664__A1 _1556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4467__A2 _0290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5011_ _0847_ _0849_ _0851_ _0852_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_97_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5416__A1 _1296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6613__B1 _2599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5913_ _1241_ _0562_ _1844_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5844_ _1754_ _1767_ _1768_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5719__A2 _0114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6767__I1 _3032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5775_ _1606_ _1628_ _1692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4726_ _0271_ _0274_ _0550_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4657_ _0342_ _3174_ _0481_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6144__A2 _1864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3608_ _2761_ _2764_ _2767_ _2768_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
X_4588_ _3101_ _0411_ _0412_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6327_ _2142_ _2139_ _2296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3539_ _2190_ _2201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3790__I _1598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5104__B1 _2922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6258_ _2219_ _2220_ _2221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5655__A1 _0287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5209_ _1068_ _3035_ _1069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_57_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6189_ _3290_ _2145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5407__A1 _0286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6080__A1 _1985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6383__A2 _2257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4394__A1 _0148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4146__A1 _2863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5894__A1 _1559_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4796__I B\[0\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4449__A2 _2763_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5646__A1 _1546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6694__I0 _2671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4082__B1 _2941_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3890_ _3047_ _3048_ _3050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4385__A1 A\[1\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5560_ _1451_ _1453_ _1456_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4511_ _0326_ _3015_ _0331_ _0333_ _0335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5491_ _0833_ _1380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4442_ _3392_ _2332_ _0266_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4373_ _0135_ _0139_ _0196_ _0197_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6112_ _1562_ _2061_ _2062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5637__A1 _0230_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6043_ _1219_ _1260_ _1986_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6062__A1 _2005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6601__A3 _2584_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6876_ _0059_ net11 net1 B\[3\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5827_ _1726_ _1748_ _1749_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_10_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3785__I _1620_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6161__I _0824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6872__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5758_ _1670_ _1671_ _1673_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4709_ _0261_ _0297_ _0533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5689_ _1595_ _0318_ _3368_ _1596_ _1597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_2_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3887__B1 _3042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5628__A1 _1470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4851__A2 _2910_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6053__A1 _1243_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5800__A1 _1716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6356__A2 _2222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4382__A4 _0960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3590__A2 _2102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5867__A1 _1765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6292__A1 _1987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5150__I _0687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4991_ _0829_ _0830_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6595__A2 _0459_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6730_ _2691_ _2698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3942_ _3035_ _3102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6661_ net8 _2645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3873_ _2299_ _3033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5612_ _1509_ _1512_ _1513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4358__A1 _0126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6592_ _1747_ _1799_ _2578_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_30_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5543_ _0070_ _1437_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5474_ _3299_ _0600_ _1361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5858__A1 _1761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4425_ _0197_ _0213_ _0249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4356_ _3372_ _0178_ _0179_ _0180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_98_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4287_ A\[0\]\[4\] _0111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6283__A1 _2007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6026_ _3252_ _3254_ _1967_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4833__A2 _0599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4597__A1 _3007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6859_ _0042_ net11 net1 B\[1\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_11_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6338__A2 _2306_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5010__A2 _0706_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3572__A2 _2545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5849__A1 _1772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6510__A2 _2427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6649__I0 _0350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5077__A2 _0922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6274__A1 _2115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4588__A1 _3101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4760__A1 _3295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3563__A2 _2419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5145__I _0628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4210_ _2921_ _3369_ _3370_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5190_ _0652_ _2984_ _1049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4141_ A\[1\]\[1\] _3301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6265__A1 _2027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4072_ _2907_ _3116_ _3232_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6017__A1 _1955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6704__I _2680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4579__A1 _3015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4974_ _0760_ _0780_ _0811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5240__A2 _1102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6713_ _2686_ _0020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3925_ _0894_ _3080_ _2987_ _3085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_32_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6644_ _2629_ _2630_ _2631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_20_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3856_ _3005_ _3015_ _3011_ _3013_ _3016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6575_ _1793_ _1783_ _2561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_30_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3787_ _2860_ _2946_ _2947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4346__A4 _2697_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3554__A2 _2354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5526_ _1318_ _1321_ _1417_ _1418_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4751__A1 _0559_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5457_ _1308_ _1337_ _1297_ _1342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_133_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4408_ _2332_ _3379_ _0232_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5388_ _3296_ _0583_ _0585_ _1265_ _1266_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_132_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4339_ _0148_ _0160_ _0162_ _0163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_59_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4806__A2 _0629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6009_ _3275_ _1947_ _1948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6815__S _2751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3490__A1 _1488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5231__A2 _1053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4034__A3 _3136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4742__A1 _0560_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6495__A1 _2437_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6247__A1 _1900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3710_ _2866_ _2869_ _2870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_18_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3784__A2 _2943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4690_ _0511_ _0513_ _0514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_119_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3641_ _2616_ _2757_ _2801_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3883__I _2070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6360_ _2327_ _2328_ _2331_ _2333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4733__A1 _0545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3572_ _2473_ _2545_ _2555_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_143_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5311_ _1116_ _1181_ _1182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_53_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6291_ _2231_ _2235_ _2257_ _2258_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_114_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6486__A1 _2467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5289__A2 _3024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5242_ _1058_ _1104_ _1105_ _1106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5173_ _0992_ _1024_ _1027_ _1028_ _1029_ _1030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_96_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4124_ _3241_ _3283_ _3284_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_111_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput1 clk net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XFILLER_84_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4055_ _3070_ _3210_ _3214_ _3215_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_37_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3472__A1 _0861_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5213__A2 _3106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4957_ _0787_ _0791_ _0792_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_71_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3908_ _3027_ _3066_ _3067_ _3068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4888_ B\[0\]\[0\] _0716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3839_ _2948_ _2998_ _1807_ _2995_ _2999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6627_ _1659_ _1660_ _2613_ _2614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_6558_ _1166_ _2542_ _2044_ _1167_ _2543_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_134_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5509_ _1395_ _1398_ _1399_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6489_ _2415_ _2412_ _2472_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4129__I net15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5452__A2 _3379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6401__A1 _2002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4007__A3 _3157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3766__A2 _2898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4799__I _0622_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4715__A1 _0285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6468__A1 _2391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6640__A1 _2500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5443__A2 _1326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3454__A1 _1169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5860_ _1778_ _1779_ _1786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4811_ B\[0\]\[6\] _0635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5791_ _1650_ _1707_ _1710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_61_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4954__A1 _0733_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4742_ _0560_ _0563_ _0565_ _0566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3757__A2 _2860_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4673_ _0495_ _0496_ _0497_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6412_ _2151_ _2388_ _2389_ _2390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4502__I _0325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3624_ _1345_ _0949_ _2784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6343_ _2311_ _2313_ _2314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3555_ _2277_ _2321_ _2365_ _2376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_143_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6274_ _2115_ _1239_ _2239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3486_ B\[3\]\[5\] _1620_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5225_ _1011_ _1012_ _1087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6829__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5682__A2 _0953_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5156_ _1003_ _1006_ _1008_ _1010_ _1011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_111_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4107_ _2959_ _3266_ _3267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5087_ _0910_ _0932_ _0934_ _0935_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4038_ _3194_ _3197_ _3198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3445__A1 _1147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3788__I _0773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6164__I _1486_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5198__A1 _1046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5989_ _1876_ _1921_ _1925_ _1926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3920__A2 _0960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5122__A1 _0886_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3987__A2 _3146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3739__A2 _2898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4164__A2 _2651_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5361__A1 _0846_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3911__A2 _2939_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5113__A1 _0963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5113__B2 _0959_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ _2893_ _0706_ _0851_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5664__A2 _1559_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6613__A1 _2597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5416__A2 _3390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6613__B2 _2491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5912_ _1482_ _1000_ _1843_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3978__A2 _3136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5843_ _1156_ _0190_ _1753_ _1767_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5774_ _1605_ _1689_ _1690_ _1691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4725_ _2930_ _3245_ _0547_ _0548_ _0549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5328__I _1199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4656_ _0472_ _0473_ _0475_ _0479_ _0480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_135_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3607_ _2766_ A\[2\]\[0\] _1180_ _1290_ _2767_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_4587_ _0152_ _0411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3538_ A\[2\]\[3\] _2190_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3902__A2 _3026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6326_ _2095_ _2097_ _2294_ _2295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5104__A1 _0953_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6257_ _1879_ _1917_ _2220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5104__B2 _0948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3469_ _1213_ _1279_ _1411_ _1422_ _1433_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_5208_ _0917_ _1068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_76_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5655__A2 _0830_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6188_ _2141_ _2143_ _2144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5139_ _0910_ _0932_ _0992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5407__A2 _0615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4918__A1 _2157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5591__A1 _0613_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5894__A2 _1569_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4449__A3 _3390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5646__A2 _1548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6694__I1 _2131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3657__A1 _2808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6733__S _2698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4909__A1 _0714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5582__A1 _0561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4385__A2 _0916_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4510_ _0332_ _0333_ _0334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_129_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5490_ _0643_ _0307_ _1379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4441_ _0079_ _2299_ _0265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4372_ _0131_ _0140_ _0196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6111_ _1897_ _1229_ _2061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5637__A2 _0706_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6042_ _1211_ _1215_ _1984_ _1985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6707__I _2678_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3663__A4 _2398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4227__I _3380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6062__A2 _1955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6875_ _0058_ net11 net1 B\[3\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5826_ _1737_ _1738_ _1748_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5757_ _1670_ _1671_ _1672_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4708_ _0250_ _0253_ _0531_ _0532_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5688_ _0958_ _1596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4639_ _0406_ _0408_ _0463_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6522__B1 _1772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3887__A1 _3038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6309_ _2273_ _2274_ _2275_ _2276_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3639__A1 _2779_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5800__A2 _1718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4119__A2 _3278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6513__B1 _2490_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3878__A1 _3037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6728__S _2692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4055__A1 _3070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4990_ _0599_ _0829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3941_ _3045_ _3101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3802__A1 _2893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6660_ _2643_ _0004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3872_ _2961_ _3032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5611_ _1508_ _1511_ _1512_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5555__A1 _1370_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4358__A2 _0141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6591_ _2268_ _2563_ _2577_ net30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5542_ _1275_ _1434_ _1435_ _1287_ _1436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_9_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5473_ _0652_ _3308_ _3305_ _0769_ _1360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4424_ _0193_ _0240_ _0247_ _0248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4355_ _0121_ _0177_ _0179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_141_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4286_ _0105_ _0109_ _0110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_58_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6025_ _2946_ _3253_ _1966_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6035__A2 _3285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4046__A1 _3202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4597__A2 _0420_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5794__B2 _1712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6858_ _0041_ net11 net1 B\[1\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_120_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5546__A1 _1247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5809_ _1630_ _1728_ _1684_ _1729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_6789_ _2731_ _2738_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_13_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5849__A2 _3369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6649__I1 _2634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6274__A2 _1239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4588__A2 _0411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5537__A1 _1427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4140_ _3299_ _0751_ _3300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6265__A2 _2030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4071_ _3229_ _3230_ _3231_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6862__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6017__A2 _1898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5776__A1 _1634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4579__A2 _0257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4973_ _0677_ _0808_ _0809_ _0810_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6712_ _2665_ _3272_ _2682_ _2686_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3924_ _3080_ _3082_ _3083_ _3071_ _3084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_60_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6643_ net14 net13 _2630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3855_ _3007_ _3015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6574_ _2556_ _2557_ _2559_ _2560_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3786_ _2945_ _2785_ _2946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4200__A1 _2945_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5525_ _1314_ _1317_ _1417_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5456_ _1337_ _1338_ _1339_ _1340_ _1341_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_59_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4407_ _0230_ _2894_ _0103_ _0231_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5387_ _1196_ _1264_ _1265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_120_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4338_ _2343_ _0161_ _0162_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6256__A2 _1915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4269_ B\[1\]\[6\] _2765_ A\[0\]\[0\] A\[0\]\[1\] _0093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_59_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4267__A1 _3324_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6008_ _3267_ _1946_ _1947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_67_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6008__A2 _1946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3490__A2 _1554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5767__A1 _1068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5519__A1 _1374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5455__B1 _0112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4325__I _3382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3640_ _2616_ _2757_ _2800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3571_ _2408_ _2505_ _2535_ _2545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_127_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5310_ _1119_ _1120_ _1181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_142_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6290_ _2251_ _2255_ _2257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_115_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5241_ _1093_ _1102_ _1105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5172_ _0909_ _1025_ _1024_ _1029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_123_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4123_ _3257_ _3282_ _3283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6238__A2 _2198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput2 execute net2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4054_ _3211_ _3213_ _3214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_56_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6715__I _2687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3472__A2 _0993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4956_ _0788_ _0789_ _0790_ _0791_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4421__A1 _0183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3907_ _3064_ _3065_ _3067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4972__A2 _0807_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4887_ _2146_ _0689_ _0715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6174__A1 _2061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6626_ _1803_ _2590_ _2613_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3838_ _2994_ _2998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6557_ _1137_ _1151_ _2542_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5921__A1 _1480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3769_ _2862_ _2870_ _2928_ _2929_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5508_ _1396_ _1397_ _1398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_106_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6488_ _2417_ _2420_ _2454_ _2471_ _2266_ net23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_10_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5439_ _1318_ _1321_ _1322_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_126_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output22_I net22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6401__A2 _1877_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4145__I A\[1\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5912__A1 _1482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4715__A2 _0295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3923__B1 _2988_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6468__A2 _2394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6712__I0 _2665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6640__A2 _2618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3454__A2 _1202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4651__A1 _0463_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6880__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4810_ B\[0\]\[6\] _0633_ A\[2\]\[0\] _1180_ _0634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_61_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5790_ _1650_ _1707_ _1709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4741_ _0265_ _0564_ _0565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4954__A2 _2004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4672_ _0482_ _0484_ _0496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_135_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6411_ _2152_ _2153_ _2177_ _2389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5903__A1 _1548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3623_ _2780_ _2782_ _2783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_128_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6342_ _2114_ _1887_ _2312_ _2200_ _2313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_3554_ _2343_ _2354_ _2365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6703__I0 _2652_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6273_ _1243_ _1996_ _2238_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3485_ _0872_ _1598_ _1609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5224_ _0974_ _1001_ _1086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5131__A2 _0873_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5155_ _1009_ _3040_ _3247_ _1005_ _1010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6646__S _2632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4890__A1 _0711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3693__A2 _2835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4106_ _3260_ _1235_ _3266_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_84_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5086_ _0929_ _0933_ _0931_ _0934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4037_ _3166_ _3195_ _3196_ _3197_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3445__A2 _1158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6871__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6395__A1 _2173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5988_ _1924_ _1925_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4939_ _2937_ _2785_ _0769_ _0770_ _0772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_21_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6609_ _2593_ _2453_ _2594_ _2595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_126_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5122__A2 _0973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3684__A2 _2843_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6862__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6310__A1 _1845_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5113__A2 _2998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5664__A3 _1569_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3675__A2 _2834_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4624__A1 _0439_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5911_ _1544_ _1551_ _1841_ _1842_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6853__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5842_ _1754_ _1755_ _1751_ _1766_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__6377__A1 _2120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5773_ _1687_ _1688_ _1690_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4724_ _3383_ _0548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4655_ _0412_ _0477_ _0478_ _0479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_3606_ _2765_ _2766_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4586_ _3043_ _3385_ _0410_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6325_ _2094_ _2141_ _2294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3537_ _2157_ _2168_ _2179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6256_ _1881_ _1915_ _2219_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3468_ _1334_ _1400_ _1422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_88_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5207_ _1006_ _1066_ _1065_ _1067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__5655__A3 _1401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6187_ _2094_ _2098_ _2142_ _2143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3666__A2 _2484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5138_ _0989_ _0990_ _0987_ _0991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_84_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6604__A2 _1801_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5069_ _0682_ _2081_ _0915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6844__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4918__A2 B\[0\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5040__A1 _0880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5591__A2 _1222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4449__A4 _0111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5646__A3 _1549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3657__A2 _2816_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3502__I _1576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4606__A1 _0419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6835__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6359__A1 _2188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5429__I _3392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6819__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5582__A2 _0972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4440_ _0165_ _0166_ _0231_ _0234_ _0264_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6531__B2 _1925_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4371_ _0142_ _0176_ _0194_ _0195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6110_ _1595_ _2058_ _2005_ _1564_ _2060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_125_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5098__A1 _0946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6041_ _1526_ _1208_ _1216_ _1984_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_6_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6598__A1 _3206_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6826__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5270__A1 _1124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6874_ _0057_ net11 net1 B\[3\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5825_ _1715_ _1746_ _1747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_22_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5022__A1 _0843_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5756_ _1359_ _1666_ _1591_ _1671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__3584__A1 _2651_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4707_ _2909_ _0530_ _0254_ _0531_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_124_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5687_ _0963_ _1595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6522__A1 _1731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4638_ _0386_ _0461_ _0462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6522__B2 _0491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4569_ _0392_ _0971_ _0393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6308_ _1526_ _2273_ _2275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6239_ _3245_ _2200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6817__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3811__A2 _2970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6513__A1 _2147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6513__B2 _2491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3878__A2 _2806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6808__I _2744_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6744__S _2706_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3940_ _3041_ _3099_ _3097_ _3100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_91_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3802__A2 _2961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3871_ _3011_ _3030_ _3031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5610_ _3351_ _0951_ _1511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6590_ _2568_ _2575_ _2546_ _2577_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4998__I _0588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5541_ _1288_ _1289_ _1435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_76_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6504__A1 _2468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5472_ _0651_ _3317_ _1359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4423_ _0195_ _0239_ _0247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_144_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3407__I B\[3\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4354_ _0121_ _0177_ _0178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_141_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4285_ _0103_ _0106_ _0108_ _0109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_101_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6024_ _3242_ _3256_ _1964_ _1965_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4294__A2 _0101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6857_ _0040_ net11 net1 B\[1\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5808_ _0282_ _1064_ _1728_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5546__A2 _0546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6788_ _2737_ _0051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5739_ _1387_ _1648_ _1652_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_136_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5537__A2 _1428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3720__A1 _2879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4070_ _2925_ _2977_ _3230_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5473__A1 _0652_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5473__B2 _0769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4972_ _0758_ _0807_ _0809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_45_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5776__A2 _1635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6711_ _2685_ _0019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3787__A1 _2860_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3923_ _2989_ _2985_ _2988_ _3081_ _3083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6642_ net2 net12 _2629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5528__A2 _0168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3854_ _3012_ _3013_ _3014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6573_ _1172_ _2558_ _2418_ _2559_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3785_ _1620_ _2945_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4200__A2 _3317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5524_ _1293_ _1324_ _1415_ _1416_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5455_ _1002_ _0161_ _0112_ _0699_ _1340_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6649__S _2632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4406_ _0229_ _0230_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5386_ _1198_ _1263_ _1264_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4337_ A\[0\]\[3\] _0161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4268_ A\[1\]\[7\] B\[3\]\[0\] _0092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6007_ _1944_ _1945_ _1946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_101_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4199_ _3322_ _3357_ _3358_ _3359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5216__A1 _0973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3600__I A\[3\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5767__A2 _0411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5519__A2 _1377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4431__I _3308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5455__A1 _1002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5455__B2 _0699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4430__A2 _0253_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4194__A1 _2939_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3570_ _2525_ _1971_ _2535_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5881__B _1581_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5240_ _1093_ _1102_ _1104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5171_ _0989_ _0990_ _1028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_116_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4122_ _3259_ _3281_ _3282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_111_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5446__A1 _1328_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4053_ _3148_ _3208_ _3212_ _3213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xinput3 input_val[0] net3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4955_ _0635_ _0734_ _2288_ _2267_ _0790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_80_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4421__A2 _0187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3906_ _3064_ _3065_ _3066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4886_ _0710_ _0711_ _0713_ _0698_ _0714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_138_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6625_ _3296_ _2608_ _2611_ _2612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3837_ _0784_ _2996_ _2997_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5347__I _0734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4251__I _3393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6556_ _1981_ _2540_ _2541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3768_ _2866_ _2869_ _2928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5507_ _0836_ _3309_ _3313_ _0837_ _1397_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_3_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6487_ _1271_ _2470_ _3296_ _2471_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3699_ _1565_ _1070_ _2859_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5438_ _1280_ _1319_ _1320_ _1321_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_134_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5685__A1 _1372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5369_ _1240_ _1242_ _1244_ _1245_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_43_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5810__I _1068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3999__A1 _3100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6641__I net3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4963__A3 _0798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6852__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5912__A2 _1000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3923__B2 _3081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5676__A1 _1528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5600__A1 _1439_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4740_ _0230_ _1235_ _0564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4671_ _0388_ _0493_ _0494_ _0495_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4167__A1 _3324_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6410_ _2152_ _2153_ _2177_ _2388_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3622_ _2781_ _1708_ _2782_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6341_ _1887_ _2281_ _2312_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3553_ A\[2\]\[1\] _2354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6500__B _2483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6272_ _1990_ _1997_ _2236_ _2237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3484_ B\[3\]\[4\] _1598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6703__I1 _3102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5667__A1 _1498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5223_ _0973_ _1083_ _1084_ _1085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5154_ _0712_ _1009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4105_ _3262_ _3264_ _3265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6873__D _0056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5085_ _0913_ _0928_ _0933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_116_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4036_ _3155_ _3165_ _3196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4642__A2 _0465_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4246__I _0069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6662__S _2638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5987_ _1923_ _1271_ _1924_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6875__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4938_ _2937_ _0769_ _0770_ _1356_ _0771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6147__A2 _2099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4869_ _2452_ _0687_ _0694_ _2092_ _0695_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_138_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4158__A1 _3317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6608_ _3210_ _3214_ _2594_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6539_ _1165_ _2521_ _2523_ _2524_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5658__A1 _1505_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4330__A1 _3274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4881__A2 _0705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5830__A1 _1729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_102_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4397__A1 _2879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5649__A1 _1536_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6697__I0 _2673_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4624__A2 _0440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5910_ _1537_ _1542_ _1841_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_34_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5841_ _1726_ _1748_ _1758_ _1765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_34_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5772_ _1687_ _1688_ _1689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4723_ _0546_ _0547_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4654_ _0408_ _0478_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3605_ B\[1\]\[7\] _2765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4585_ _0406_ _0408_ _0409_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6324_ _2287_ _2292_ _2293_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3536_ B\[1\]\[0\] _2168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4560__A1 _3297_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6688__I0 _2665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6255_ _2191_ _2194_ _2217_ _2218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_89_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3467_ _1334_ _1400_ _1411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5206_ _3008_ _0800_ _1066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6186_ _2090_ _2091_ _2089_ _2142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5137_ _0675_ _3025_ _0990_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6065__A1 _2001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5068_ _0889_ _0890_ _0914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_input14_I sel_in[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5812__A1 _1729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4019_ _3173_ _3178_ _3179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5591__A3 _0354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4303__A1 _3251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6056__A1 _0857_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5803__A1 _0387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4606__A2 _0428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5031__A2 _0873_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4790__A1 _0613_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4542__A1 _0363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4370_ _0145_ _0175_ _0194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5098__A2 _0982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6295__A1 _2258_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6040_ _1935_ _1979_ _1981_ _1983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I input_val[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5270__A2 _1135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6873_ _0056_ net11 net1 B\[3\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5824_ _1725_ _1744_ _1745_ _1746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_50_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5755_ _1666_ _1667_ _1668_ _1669_ _1670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_72_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3584__A2 _2660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4706_ _0257_ _0530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5686_ _1592_ _1593_ _1594_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4637_ _0389_ _0461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6522__A2 _0490_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4568_ A\[1\]\[2\] _0392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3519_ _1971_ _1982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6307_ _2058_ _0670_ _2274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_103_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4499_ _0321_ _0322_ _0323_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6286__A1 _1200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5089__A2 _0936_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6238_ _2114_ _2198_ _2199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6169_ _2116_ _2122_ _2123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6038__A1 _1935_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5013__A2 _0798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6210__A1 _1957_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3575__A2 _2565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6513__A2 _2485_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4524__A1 _0325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5721__B1 _0149_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6277__A1 _2115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6096__I _2043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6029__A1 _0979_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5252__A2 _1112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3870_ _3004_ _3006_ _3030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5004__A2 _0802_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6201__A1 _1239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5540_ _1248_ _0281_ _1434_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4763__A1 _0586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5471_ _0649_ A\[1\]\[4\] _1358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4422_ _0188_ _0192_ _0245_ _0246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4353_ _0142_ _0176_ _0177_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4284_ _0107_ _1971_ _0108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6023_ _3250_ _3255_ _1964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_100_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3423__I _0916_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4294__A3 _0117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6815__I0 _1877_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6440__A1 _2414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6856_ _0039_ net11 net1 B\[0\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_22_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5807_ _0980_ _0257_ _1727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6787_ _0830_ _2640_ _2733_ _2737_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3999_ _3100_ _3158_ _3159_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5738_ _1650_ _1651_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5669_ _1503_ _1506_ _1575_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4506__A1 _3326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6259__A1 _2218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3493__A1 _1136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6806__I0 _2940_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3796__A2 _2896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4993__A1 _0643_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3720__A2 _2288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5473__A2 _3308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6422__A1 _2268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5225__A2 _1012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4971_ _0758_ _0807_ _0808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_91_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6710_ _2663_ _3247_ _2682_ _2685_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_63_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3787__A2 _2946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4984__A1 _0774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3922_ _3081_ _2989_ _3082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3853_ _0806_ _1114_ _3013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6641_ net3 _2628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5528__A3 _1310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6572_ _1167_ _1171_ _2368_ _2558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3784_ _2942_ _2943_ _2944_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5523_ _1307_ _1322_ _1415_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6489__A1 _2415_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5454_ _3323_ _0690_ _1339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4405_ _0164_ _0229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5385_ _1204_ _1207_ _1262_ _1263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_132_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4336_ _3392_ _2644_ _0160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4249__I _0072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6665__S _2631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4267_ _3324_ _0089_ _0090_ _0066_ _0091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6110__B1 _2005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6006_ _3263_ _3274_ _1945_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4198_ _3338_ _3356_ _3358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4975__A1 _0764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6839_ _0022_ net11 net1 A\[2\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4727__A1 _0549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3950__A2 _3107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5543__I _0070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5455__A2 _0161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3466__A1 _1378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4194__A2 _3353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5694__A2 _1602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5170_ _0909_ _1025_ _1027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4121_ _3268_ _3280_ _3281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_110_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6643__A1 net14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4052_ _3151_ _3152_ _3212_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_111_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 input_val[1] net4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4954_ _0733_ _2004_ _0789_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3905_ _1851_ _2837_ _3065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4885_ _2525_ _0686_ _0712_ _2452_ _0713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_71_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6624_ _2225_ _2610_ _2611_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3836_ _2994_ _2995_ _2996_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5382__A1 _1236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6555_ _2529_ _2539_ _2540_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3767_ _2873_ _2899_ _2926_ _2927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5506_ _1380_ _0255_ _0128_ _0870_ _1396_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_106_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6486_ _2467_ _2469_ _2470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3698_ _2804_ _2856_ _2857_ _2858_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5134__A1 _0983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5437_ _0997_ _3387_ _1320_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5363__I _2893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5368_ _0847_ _1243_ _1244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3696__A1 _2808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4319_ _0101_ _0117_ _0143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5299_ _1124_ _1135_ _1168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6634__A1 _0304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5437__A2 _3387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3448__A1 _1180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3767__B _2926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3620__A1 _0707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3923__A2 _2985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5273__I _1064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6625__A1 _3296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3439__A1 _1059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3521__I _1993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5600__A2 _1442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3611__A1 _2759_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4670_ _0489_ _0492_ _0494_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3621_ _1532_ _1598_ _2781_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5364__A1 _1239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4167__A2 _3326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3552_ _2332_ _2343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6340_ _0564_ _1890_ _2204_ _2205_ _2209_ _2311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_116_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6271_ _1998_ _2010_ _2236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3483_ _1565_ _1576_ _1587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5222_ _1075_ _1076_ _1084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5153_ _3106_ _1007_ _1008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6616__A1 _3070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5419__A2 B\[0\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4104_ _3263_ _3264_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5084_ _0930_ _0931_ _0932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_111_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4035_ _3167_ _3179_ _3195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4527__I _0328_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3431__I _1004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3850__A1 _1202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5986_ net16 _1923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4937_ _0649_ _0770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4868_ _0693_ _0694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6607_ _3210_ _3214_ _2593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5355__A1 _1229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4158__A2 _0927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3819_ _2914_ _2978_ _2979_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4799_ _0622_ _0623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6538_ _3191_ _2522_ _1273_ _2523_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6189__I _3290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5107__A1 _0955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6469_ _2448_ _2450_ _2451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_133_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5658__A2 _1562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3669__A1 _2387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4330__A2 _2809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4881__A3 _0708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4094__A1 _2946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5830__A2 _1732_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3841__A1 _2991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6652__I _2631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4397__A2 _0220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3516__I A\[2\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6763__S _2719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5821__A2 _1699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5840_ _1715_ _1746_ _1764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_62_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5585__A1 _1482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5771_ _1338_ _1682_ _1632_ _1688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_99_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4722_ _0220_ _0546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4653_ _0476_ _3169_ _0477_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3604_ _2762_ _2763_ A\[2\]\[0\] A\[2\]\[1\] _2764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4584_ _0351_ _0407_ _0350_ _3169_ _0408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__3899__A1 _3029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6323_ _2106_ _2290_ _2291_ _2292_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3535_ _2146_ _2157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4560__A2 _2940_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3426__I _0949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6688__I1 _1817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3466_ _1378_ _1389_ _1400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6254_ _2211_ _2216_ _2217_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_88_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5205_ _1064_ _2932_ _1065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_130_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6185_ _2139_ _2140_ _2141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5136_ _0987_ _0988_ _0989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5067_ _0911_ _0912_ _0913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_38_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4076__A1 _2936_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6842__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5812__A2 _1732_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4018_ _3176_ _3177_ _3178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5576__A1 _1418_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5969_ _1892_ _1903_ _1904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_32_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5591__A4 _0357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4000__A1 _3093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4303__A2 _3311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5500__A1 _1293_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5803__A2 _1596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5567__A1 _1394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5319__A1 _0907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4542__A2 _0364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6865__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4058__B2 _3211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6598__A3 _2582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6872_ _0055_ net11 net1 B\[2\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__5558__A1 _1381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5823_ _1742_ _1743_ _1745_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5754_ _3297_ _0830_ _1669_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4705_ _0246_ _0300_ _0528_ _0529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_136_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5685_ _1372_ _1588_ _1361_ _1593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_120_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4636_ _0419_ _0428_ _0402_ _0460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_135_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4567_ _0387_ _0319_ _0391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6306_ _2126_ _2127_ _2061_ _2273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3518_ B\[1\]\[0\] _1971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4498_ _0310_ _0311_ _0322_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6286__A2 _2003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6237_ _3243_ _2198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5371__I _0731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3449_ _1169_ _1202_ _1213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_76_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6168_ _2117_ _2118_ _2121_ _2122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5119_ _0969_ _0970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4049__A1 _3148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6099_ _1811_ _1817_ _1825_ _2047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_17_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5797__A1 _0314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5549__A1 _1439_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4221__A1 _3037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5721__A1 _0694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4524__A2 _3007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5721__B2 _0687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6277__A2 _2160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6029__A2 _2908_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4460__A1 _0219_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6201__A2 _3243_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4763__A2 _1796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5470_ _1352_ _1355_ _1357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_129_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4421_ _0183_ _0187_ _0245_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_99_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4352_ _0145_ _0175_ _0176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_140_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4283_ A\[0\]\[7\] _0107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4279__A1 _0102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6022_ _1942_ _1962_ _1963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_100_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6815__I1 _2649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5779__A1 _1691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6440__A2 _2416_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6855_ _0038_ net11 net1 B\[0\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6750__I _2705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5806_ _1721_ _1724_ _1726_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6786_ _2736_ _0050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3998_ _3097_ _3103_ _3158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5737_ _1618_ _1621_ _1650_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_129_36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5668_ _1504_ _1505_ _1574_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4619_ _0431_ _0441_ _0443_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5703__A1 _1612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6751__I0 _2665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5599_ _1399_ _1408_ _1497_ _1498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6806__I1 _2640_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4442__A1 _3392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4993__A2 _2943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6660__I _2643_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4745__A2 _0568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6742__I0 _2652_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5170__A2 _1025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6422__A2 _2301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4970_ _0781_ _0805_ _0807_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_91_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3921_ _1576_ _3081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6640_ _2500_ _2618_ _2620_ _2626_ _1269_ net18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3852_ _3005_ _3007_ _3011_ _3012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5528__A4 _1002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6571_ _0506_ _2226_ _2557_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4736__A2 _3033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5933__A1 _1864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3783_ _1532_ _2943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5522_ _1394_ _1409_ _1413_ _1414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_30_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5453_ _1310_ _0088_ _1338_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6733__I0 _2669_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4404_ _0163_ _0172_ _0227_ _0228_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5384_ _1217_ _1261_ _1262_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4335_ _0110_ _0116_ _0158_ _0159_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3434__I A\[3\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6110__A1 _1595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4266_ _0064_ _0067_ _0090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6110__B2 _1564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6745__I _2708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6005_ _3269_ _3244_ _1944_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4197_ _3338_ _3356_ _3357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4672__A1 _0482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6681__S _2656_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4975__A2 _0779_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6838_ _0021_ net11 net1 A\[2\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__6177__A1 _2131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5924__A1 _1847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6769_ _2717_ _2724_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_10_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6724__I0 _2658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6655__I net6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3466__A2 _1389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5207__A3 _1065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6168__A1 _2117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5915__A1 _1539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3519__I _1971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6340__A1 _0564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4120_ _2970_ _3279_ _3280_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_110_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6643__A2 net13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4051_ _3027_ _3066_ _3211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_110_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput5 input_val[2] net5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4085__I _3244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4953_ _0731_ _2026_ _0788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3904_ _3028_ _3059_ _3061_ _3062_ _3063_ _3064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__6159__A1 _1845_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4884_ _0692_ _0712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6623_ _1036_ _2609_ _2610_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5906__A1 _0287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3835_ _2950_ _2995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3429__I _0828_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6554_ _3166_ _3195_ _2539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3766_ _2875_ _2898_ _2926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5505_ _1228_ _3311_ _1395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6485_ _2323_ _2333_ _2468_ _2469_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3697_ _2808_ _2816_ _2857_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5436_ _0848_ _0220_ _1319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5134__A2 _0986_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5367_ _0888_ _3260_ _1243_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3696__A2 _2816_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4893__A1 _0704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4318_ _0124_ _0126_ _0141_ _0142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_5298_ _1137_ _1166_ _1167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6634__A2 _0525_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4249_ _0072_ _0073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3448__A2 _1191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6874__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4723__I _0546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3620__A2 _0905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6625__A2 _2608_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4636__A1 _0419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6865__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3620_ _0707_ _0905_ _2780_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5364__A2 _0999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3693__B _2852_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4572__B1 _3072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3551_ B\[1\]\[5\] _2332_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6270_ _2232_ _2233_ _2235_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3482_ A\[3\]\[1\] _1576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5221_ _1075_ _1076_ _1083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4875__A1 _0697_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3678__A2 _2836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5152_ _0800_ _1007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4103_ _2821_ _3263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5083_ _0704_ _0721_ _0679_ _0931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_57_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4034_ _3090_ _3127_ _3136_ _3194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_37_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6856__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3850__A2 _3009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5985_ _1876_ _1921_ _1922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_52_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5052__A1 _0893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4936_ _0655_ _0769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4867_ _0692_ _0693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6606_ _2590_ _2591_ _2592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3818_ _2925_ _2977_ _2978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5355__A2 _3004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4798_ B\[0\]\[5\] _0622_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6537_ _3189_ _3190_ _2145_ _2522_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3749_ _2908_ _2909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6304__A1 _2111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5107__A2 _0956_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6468_ _2391_ _2394_ _2449_ _2450_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5419_ A\[0\]\[6\] B\[0\]\[0\] _1300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6399_ _2165_ _2166_ _1957_ _2375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3669__A2 B\[1\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4330__A3 _0152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6847__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4094__A2 _3253_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3841__A2 _2992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output20_I net20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5043__A1 _0621_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5594__A2 _1492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6838__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3832__A2 _2982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5034__A1 _0905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5770_ _1682_ _1683_ _1684_ _1685_ _1687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_62_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5585__A2 _1007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3596__A1 _2718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4721_ _0208_ _0209_ _0288_ _0294_ _0545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_30_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4652_ _0351_ _0476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3603_ B\[1\]\[7\] _2763_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4583_ _3101_ _0407_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3899__A2 _3057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6322_ _2289_ _2137_ _2291_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3534_ A\[2\]\[5\] _2146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6253_ _2213_ _2215_ _2216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3465_ B\[3\]\[0\] _1389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4848__A1 _0670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5204_ _1009_ _1064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6184_ _2104_ _2105_ _2138_ _2140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5135_ _0983_ _0986_ _0988_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5066_ _0617_ _0892_ _0912_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6829__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4076__A2 _2954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4017_ _3168_ _3172_ _3177_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_84_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5968_ _1896_ _1902_ _1903_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4919_ _0622_ _2201_ _0750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5899_ _1553_ _1570_ _1827_ _1828_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4000__A2 _2849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4839__A1 _0611_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3511__A1 _1422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4067__A2 _2919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5264__A1 _1062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6663__I _2646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3814__A2 _2973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5016__A1 _0635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3578__A1 _2376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6516__A1 _3186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3527__I _1938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6774__S _2724_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4058__B3 _3213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3805__A2 _2890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6871_ _0054_ net11 net1 B\[2\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5822_ _1742_ _1743_ _1744_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_35_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5753_ _0948_ _0395_ _0953_ _3367_ _1668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4704_ _0248_ _0299_ _0528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6507__A1 _2361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5684_ _1588_ _1589_ _1590_ _1591_ _1592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_136_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4635_ _0454_ _0457_ _0458_ _0459_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_116_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4566_ _0386_ _0389_ _0390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5730__A2 _1640_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6305_ _2270_ _2136_ _2271_ _2272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3517_ _1938_ _1949_ _1960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4497_ _0316_ _0320_ _0321_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6236_ _0564_ _1890_ _2197_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3448_ _1180_ _1191_ _1202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5494__A1 _1381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6684__S _2656_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6167_ _2119_ _2120_ _2121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5118_ _0615_ _0969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6098_ _1980_ _1983_ _2036_ _2045_ _2046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5246__A1 _1100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5049_ _0887_ _0891_ _0892_ _0617_ _0893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_85_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5797__A2 _0953_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5099__I _0597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5549__A2 _1442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4221__A2 _3380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5721__A2 _0220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6658__I net7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5485__A1 _1363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4420_ _3371_ _0242_ _0243_ _0244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__6832__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3723__A1 _1290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4351_ _0157_ _0174_ _0175_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4282_ _0072_ _2484_ _0106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4279__A2 _2398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5476__A1 A\[1\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6021_ _1951_ _1961_ _1962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_101_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5779__A2 _1694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6854_ _0037_ net11 net1 B\[0\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_62_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5805_ _1722_ _1724_ _1725_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6785_ _1039_ _2637_ _2733_ _2736_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5400__A1 _0149_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3997_ _3074_ _3156_ _3157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4551__I _0374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5736_ _1387_ _1648_ _1649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5951__A2 _0573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3962__A1 _3047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5667_ _1498_ _1515_ _1572_ _1573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4618_ _0431_ _0441_ _0442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5598_ _1403_ _1407_ _1497_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5703__A2 _1156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6751__I1 _1000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3714__A1 _2820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4911__B1 _0682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4549_ _3373_ _0372_ _0373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6219_ _2151_ _2154_ _2177_ _2178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_89_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3630__I A\[3\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4442__A2 _2332_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6855__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3953__A1 _3104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5155__B1 _3247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6742__I1 _1731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3705__A1 _2760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4902__B1 _2026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5458__A1 _1341_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3920_ _2984_ _0960_ _3080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3851_ _3010_ _3011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4197__A1 _3338_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6570_ _0499_ _0505_ _2556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3782_ _1565_ _2942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5933__A2 _1865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5521_ _1384_ _1410_ _1412_ _1413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3944__A1 _3097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5452_ _0692_ _3379_ _1337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6733__I1 _0979_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5697__A1 _1326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4403_ _0167_ _0171_ _0227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5383_ _1219_ _1260_ _1261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_132_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4334_ _0105_ _0109_ _0158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4265_ _0088_ _3033_ _0089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4121__A1 _3268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6004_ _3268_ _3280_ _1943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4196_ _3343_ _3349_ _3355_ _3356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_68_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6878__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6837_ _0020_ net11 net1 A\[2\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_11_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6177__A2 _0670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6768_ _2723_ _0043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5719_ _0917_ _0114_ _1630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6699_ net13 _2675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6724__I1 _1829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3625__I _1499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4360__A1 _1620_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6101__A2 _1858_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5612__A1 _1509_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6671__I net12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6168__A2 _2118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4179__A1 _0707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5915__A2 _1845_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3926__A1 _3084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3535__I _2146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4050_ _3154_ _3205_ _3207_ _3209_ _3210_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_110_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4366__I _0189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput6 input_val[3] net6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4952_ _0708_ _0785_ _0786_ _0750_ _0787_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_75_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3903_ _1862_ _3060_ _3059_ _3063_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_4883_ _2515_ _0681_ _0711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6622_ _1184_ _1186_ _2597_ _2609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3834_ A\[3\]\[0\] _2994_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5906__A2 _0959_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6553_ _0499_ _2491_ _2537_ _2538_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3765_ _2920_ _2924_ _2925_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5504_ _1277_ _1292_ _1393_ _1394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6484_ _2317_ _2322_ _2468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3696_ _2808_ _2816_ _2856_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5435_ _1314_ _1317_ _1318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_134_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6331__A2 _2300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4342__A1 _0102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5366_ _1241_ _3264_ _1242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4893__A2 _0721_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4317_ _0131_ _0140_ _0141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_43_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5297_ _1153_ _1165_ _1166_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_59_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6095__A1 _1923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4248_ A\[0\]\[5\] _0072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5842__A1 _1754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4179_ _0707_ _3301_ _3339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6440__B _2418_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4581__A1 _0282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6666__I _2648_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5833__A1 _1754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4636__A2 _0428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6615__B _2593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4939__A3 _0769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3550_ _2288_ _2310_ _2321_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4572__A1 _2983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4572__B2 _3367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3481_ B\[3\]\[6\] _1565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6313__A2 _2118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4324__A1 _0111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5220_ _0970_ _3116_ _1082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4875__A2 _0701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5151_ _1005_ _3246_ _1006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4102_ _2343_ _3262_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5082_ _0913_ _0928_ _0929_ _0930_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4033_ _3166_ _3192_ _3193_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_37_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5984_ _1918_ _1920_ _1921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4935_ _0765_ _0767_ _0768_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_36_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4866_ B\[0\]\[1\] _0692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6605_ _1714_ _1801_ _2591_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6260__B _2222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3817_ _2927_ _2976_ _2977_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4797_ _2882_ _0620_ _0621_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3748_ _2907_ _2908_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6536_ _1163_ _1164_ _2044_ _2521_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6467_ _2386_ _2390_ _2449_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3679_ _1851_ _2837_ _2838_ _2839_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_5418_ _1294_ _1295_ _1297_ _1298_ _1299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6398_ _2372_ _2373_ _2374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5349_ _1222_ _1223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5390__I _1267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4330__A4 _0114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6068__A1 _1227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4618__A2 _0441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5043__A2 _0886_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5034__A2 _0829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5585__A3 _1309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3596__A2 _2746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4793__A1 _0614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4720_ _0278_ _0296_ _0543_ _0544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4651_ _0463_ _0474_ _0475_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_3602_ B\[1\]\[6\] _2762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4582_ _0355_ _0404_ _0405_ _0406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_3533_ _1960_ _2015_ _2059_ _2124_ _2135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_6321_ _2289_ _2137_ _2290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6298__A1 _2224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6298__B2 _0585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6252_ _1896_ _1901_ _2214_ _2215_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3464_ _1367_ _1378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4848__A2 _2910_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5203_ _1062_ _2923_ _1063_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6183_ _2104_ _2105_ _2138_ _2139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5134_ _0983_ _0986_ _0987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_69_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5065_ _0887_ _0891_ _0911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3808__B1 _2430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4016_ _3082_ _3175_ _3156_ _3176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_65_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5967_ _1899_ _1901_ _1902_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4918_ _2157_ B\[0\]\[3\] _0749_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5898_ _1536_ _1552_ _1827_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4849_ _0663_ _0667_ _0672_ _0673_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6519_ _1069_ _1157_ _2504_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5264__A2 _2849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5016__A2 _0633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6516__A2 _2453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6790__S _2738_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6870_ _0053_ net11 net1 B\[2\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_90_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5007__A2 _0618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6204__A1 _3243_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5821_ _1698_ _1699_ _1679_ _1743_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_50_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5752_ _3367_ _1043_ _1667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4703_ _0304_ _0525_ _0526_ _0527_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5683_ _0307_ _0951_ _1591_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4634_ _0374_ _0376_ _0458_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5191__A1 _1042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4565_ _0385_ _0388_ _0389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_128_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6304_ _2111_ _2130_ _2271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3516_ A\[2\]\[4\] _1949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3741__A2 _2900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4496_ _0317_ _0318_ _3368_ _0319_ _0320_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3447_ B\[1\]\[4\] _1191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6235_ _1885_ _1891_ _2195_ _2196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5494__A2 _1382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6166_ _1223_ _2120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6764__I _2721_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5117_ _0957_ _0967_ _0968_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6097_ _2038_ _2042_ _2044_ _2045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6443__A1 _2337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5246__A2 _1101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5048_ _0614_ _0616_ _0892_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input12_I sel_in[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5485__A2 _1358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3496__A1 _1587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6809__I0 _0319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3799__A2 _1191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4996__A1 _0766_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6342__C _2200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3420__A1 _0861_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4350_ _0159_ _0173_ _0174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__3723__A2 _2766_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4920__A1 _0727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4281_ _3394_ _0103_ _0104_ _0078_ _0105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_98_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5476__A2 _0655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6020_ _1954_ _1959_ _1961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3487__A1 _1620_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input4_I input_val[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5228__A2 _1089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4987__A1 _0824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6853_ _0036_ net11 net1 B\[0\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_90_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4739__A1 _0562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5804_ _1723_ _1673_ _1724_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6784_ _2735_ _0049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3996_ _3077_ _3156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5735_ _1350_ _1390_ _1648_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_50_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3411__A1 _0762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3962__A2 _3048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5666_ _1502_ _1514_ _1572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_108_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4617_ _0436_ _0439_ _0440_ _0441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_135_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5597_ _1474_ _1495_ _1496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5703__A3 _1607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3714__A2 _2832_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4911__B2 _2690_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4548_ _0087_ _0118_ _0372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_132_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4479_ _0302_ _0303_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5467__A2 _0588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6218_ _2171_ _2176_ _2177_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_58_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6149_ _0685_ _2101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6416__A1 _1935_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6416__B2 _2182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_78 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3953__A2 _3112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5155__A1 _1009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4902__A1 _0731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3705__A2 _1356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4902__B2 _0612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4969__A1 _0783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3641__A1 _2616_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4652__I _0351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3850_ _1202_ _3009_ _3010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4197__A2 _3356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3781_ _2938_ _2940_ _2784_ _2941_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_13_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5520_ _1374_ _1377_ _1412_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3944__A2 _3100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5451_ _1328_ _1329_ _1336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_67_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4402_ _0154_ _0225_ _0226_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5382_ _1236_ _1259_ _1260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_126_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4333_ _0147_ _0156_ _0157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_141_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4264_ A\[0\]\[3\] _0088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6003_ _3257_ _3282_ _1941_ _1942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4827__I _0596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4195_ _3347_ _3352_ _3354_ _3355_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_67_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6836_ _0019_ net11 net1 A\[2\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6767_ _2640_ _3032_ _2719_ _2723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3979_ _3090_ _3137_ _3138_ _3139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5718_ _0693_ _3390_ _1629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6698_ _2674_ _0015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5137__A1 _0675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5649_ _1536_ _1552_ _1553_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_105_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3699__A1 _1565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4360__A2 A\[1\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6637__A1 _3221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4737__I _0168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3871__A1 _3011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6822__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5073__B1 _3271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3623__A1 _2780_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5376__A1 _0847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4179__A2 _3301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3926__A2 _3085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4351__A2 _0174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5851__A2 _1039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput7 input_val[4] net7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3862__A1 _3017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5603__A2 _0256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4951_ _0727_ _0749_ _0786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3902_ _3023_ _3026_ _3062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4882_ _2704_ _0686_ _0710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6621_ _0383_ _2607_ _2608_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5367__A1 _0888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3833_ _2991_ _2992_ _2993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6552_ _0498_ _2536_ _2537_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3764_ _2921_ _2923_ _2924_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5503_ _1286_ _1291_ _1393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4590__A2 _0412_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6483_ _2465_ _2466_ _2467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3695_ _2789_ _2793_ _2854_ _2855_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5434_ _1309_ _1315_ _1316_ _1317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_69_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4342__A2 _2037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5365_ _0888_ _1241_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6619__A1 _0514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4316_ _0135_ _0139_ _0140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_87_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5296_ _1163_ _1164_ _1165_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_141_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6095__A2 _1271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4247_ _1982_ _0070_ _0071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3461__I A\[3\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6845__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4178_ _3327_ _3331_ _3336_ _3337_ _3338_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_83_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6819_ _0002_ net11 net1 A\[0\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4030__A1 _3176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4581__A2 _3096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4869__B1 _0694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5530__A1 _0164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4939__A4 _0770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4572__A2 _0395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3480_ _1521_ _1455_ _1543_ _1554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_143_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4324__A2 _1191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6868__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3532__B1 _2092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5150_ _0687_ _1005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4101_ _3260_ _3034_ _3261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5081_ _0925_ _0926_ _0929_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_57_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4088__A1 _3243_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4032_ _3180_ _3191_ _3192_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5983_ _0532_ _0579_ _1919_ _1920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4934_ _0664_ _0766_ _0767_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_127_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4865_ _0690_ _2806_ _0691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6604_ _1714_ _1801_ _2590_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3816_ _2955_ _2975_ _2976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4012__A1 _3107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4796_ B\[0\]\[3\] _0620_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6535_ _0497_ _2491_ _2519_ _2520_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3747_ B\[3\]\[7\] _2907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4061__B _3220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6466_ _2446_ _2447_ _2448_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3678_ _2777_ _2836_ _2838_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_134_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5417_ _0073_ _0699_ _0712_ _3380_ _1298_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5512__A1 _1401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6397_ _2171_ _2176_ _2373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5348_ _1221_ _1222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5279_ _1050_ _1145_ _1126_ _1146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_47_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5815__A2 _1734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3826__A1 _2983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6240__A2 _2200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5751__A1 _0392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6677__I net4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5503__A1 _1286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4242__A1 _2343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4793__A2 _0616_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4650_ _3181_ _0189_ _0474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput10 input_val[7] net10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3601_ _2760_ _1389_ _2761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4545__A2 _0368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4581_ _0282_ _3096_ _0405_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6790__I0 _1596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6320_ _2109_ _2289_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_128_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3532_ _2070_ _2004_ _2092_ _2113_ _2124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6251_ _1899_ _2214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3463_ _1356_ _1367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5491__I _0833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5202_ _0969_ _1062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6182_ _2106_ _2109_ _2137_ _2138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_112_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5133_ _0984_ _0985_ _0986_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5064_ _0909_ _0910_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3808__A1 _2879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6536__B _2044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3808__B2 _2812_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4015_ _3025_ _3174_ _3175_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4481__A1 _0971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5966_ _0290_ _1900_ _1901_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5430__B1 _1002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4917_ _0744_ _0747_ _0748_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5897_ _1819_ _1825_ _1826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_139_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4848_ _0670_ _2910_ _0671_ _0672_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4779_ _0594_ _0828_ _0603_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6781__I0 _1772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6518_ _0490_ _0407_ _0472_ _0491_ _2503_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_4_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6449_ _2342_ _2428_ _2429_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_106_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6461__A2 _2385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4472__A1 _0280_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4224__A1 _3045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5972__A1 _0545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5724__A1 _1634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6772__I0 _2645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5660__B1 _0958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6204__A2 _2160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5820_ _1726_ _1739_ _1740_ _1742_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5751_ _0392_ _0946_ _1666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4702_ _0244_ _0301_ _0526_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5682_ _0395_ _0953_ _0256_ _1042_ _1590_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6507__A3 _2433_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5715__A1 _0325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4633_ _0446_ _0455_ _0456_ _0457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6763__I0 _2634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5191__A2 _3081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4564_ _0387_ _3075_ _0388_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6303_ _2111_ _2130_ _2270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3515_ _1927_ _1938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3734__I _2037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4495_ _2995_ _0319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6234_ _1892_ _1903_ _2195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3446_ A\[2\]\[1\] _1180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6165_ _0562_ _2119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5116_ _0965_ _0966_ _0967_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6096_ _2043_ _2044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6443__A2 _2355_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5047_ _0889_ _0890_ _0891_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4454__A1 _0263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6780__I _2731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4757__A2 _0580_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5954__A1 _1886_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5949_ _0559_ _0574_ _1882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5182__A2 _1039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6809__I1 _2642_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4996__A2 _0834_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6690__I net8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5945__A1 _1877_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3420__A2 _0883_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6370__A1 _0670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4381__B1 _0960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3723__A3 _2882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4280_ _0080_ _2419_ _3037_ _3393_ _0104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6673__A2 _2654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3487__A2 _0740_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4436__A1 _0216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4987__A2 _2933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6852_ _0035_ net11 net1 B\[0\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5803_ _0387_ _1596_ _1723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4739__A2 _3262_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6783_ _1043_ _2634_ _2733_ _2735_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3995_ _3115_ _3124_ _3091_ _3155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_22_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5734_ _1625_ _1645_ _1646_ _1647_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_50_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3411__A2 _0784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5665_ _1553_ _1570_ _1571_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5944__I _2909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4616_ _0349_ _0365_ _0440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6361__A1 _2323_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5596_ _1485_ _1494_ _1495_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_85_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4911__A2 _0716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4547_ _0347_ _0369_ _0370_ _0371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3464__I _1367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6113__A1 _2060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4478_ _0244_ _0301_ _0302_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6775__I _2728_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6217_ _2173_ _2175_ _2176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_89_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3429_ _0828_ _0993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6148_ _1929_ _2046_ _1270_ _2100_ net20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6079_ _1987_ _2024_ _2025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_57_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6015__I _2938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4902__A2 _2354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3705__A3 _1510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6407__A2 _2383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4969__A2 _0804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3641__A2 _2757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5918__A1 _1221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3549__I _2299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6591__A1 _2268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3780_ _2939_ _2940_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3944__A3 _3103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5450_ _1331_ _1333_ _1335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4401_ _0219_ _0224_ _0225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6796__S _2738_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5381_ _1238_ _1258_ _1259_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_132_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4332_ _0151_ _0155_ _0156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_125_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4263_ _3377_ _0085_ _0086_ _0087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_114_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4657__A1 _0342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6002_ _3259_ _3281_ _1941_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4194_ _2939_ _3353_ _3354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4409__A1 _0102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5082__A1 _0913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3632__A2 _0916_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6835_ _0018_ net11 net1 A\[2\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_39_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5909__A1 _1830_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3459__I _1246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6582__A1 _2564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6766_ _2722_ _0042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3978_ _3127_ _3136_ _3138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5717_ _0411_ _0998_ _1000_ _0328_ _1628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6697_ _2673_ _2058_ _2666_ _2674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5648_ _1544_ _1551_ _1552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5137__A2 _3025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4345__B1 _2697_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5579_ _1426_ _1430_ _1475_ _1476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4896__A1 _0632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3699__A2 _1070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6877__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5073__A1 _0694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6454__B _2433_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5073__B2 _0917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4820__A1 _0643_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6573__A1 _1172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5584__I _0230_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6325__A1 _2094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4887__A1 _2146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6629__B _2615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6628__A2 _2614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4639__A1 _0406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5300__A2 _1151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6868__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput8 input_val[5] net8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4950_ _2157_ B\[0\]\[4\] _0785_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3614__A2 _2773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3901_ _1862_ _3060_ _3061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4881_ _0619_ _0705_ _0708_ _0709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_33_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6620_ _2604_ _2605_ _2607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3832_ _1466_ _2982_ _0938_ _2992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_60_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5367__A2 _3260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6551_ _0470_ _0502_ _2536_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3763_ _2922_ _2923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5502_ _1325_ _1350_ _1351_ _1388_ _1391_ _1392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_6482_ _2456_ _2457_ _2464_ _2466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
X_3694_ _2783_ _2794_ _2854_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5433_ _0073_ _1296_ _1316_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4878__A1 _0622_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5364_ _1239_ _0999_ _1240_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3550__A1 _2288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4315_ _0132_ _0137_ _0138_ _0139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_114_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5295_ _1146_ _1148_ _1164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_141_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4246_ _0069_ _0070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6859__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4177_ _3332_ _3335_ _3337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5055__A1 _0587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4802__A1 _0625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6818_ _0001_ net11 net1 A\[0\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6749_ _2710_ _0035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4869__A1 _2452_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4869__B2 _2092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3541__A1 _2179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3652__I _2762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5046__A1 _0621_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4483__I _3301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3532__A1 _2070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3532__B2 _2113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3562__I _2387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4100_ _2892_ _3260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5080_ _0925_ _0926_ _0928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_97_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4088__A2 _3245_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4031_ _3189_ _3190_ _3191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_96_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5982_ _0534_ _0578_ _1919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_53_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4933_ _1444_ B\[2\]\[4\] _0766_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6537__A1 _3189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4864_ _0689_ _0690_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6603_ _2103_ _2578_ _2589_ _1270_ net31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3815_ _2957_ _2974_ _2975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4795_ _2201_ _0618_ _0619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4012__A2 _3170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6534_ _0495_ _0496_ _2519_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_20_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3746_ _2904_ _2905_ _2906_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_107_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6465_ _2442_ _2445_ _2447_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3677_ _2777_ _2836_ _2837_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_134_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5416_ _1296_ _3390_ _1297_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6396_ _2156_ _2170_ _2372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5512__A2 _1363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5347_ _0734_ _1221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5278_ _3024_ _1039_ _1145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5276__A1 _1073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4229_ _3381_ _3384_ _3386_ _3388_ _3389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3826__A2 _2985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5399__I _0627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5751__A2 _0946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6700__A1 net14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6693__I net9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3817__A2 _2976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5019__A1 _0790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4242__A2 _0065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6519__A1 _1069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6835__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3600_ A\[3\]\[7\] _2760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput11 reset net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_20
X_4580_ _0328_ _3098_ _0404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6790__I1 _2642_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3531_ _2102_ _2113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6250_ _2131_ _2172_ _2213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3462_ _1345_ _1356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5201_ _1060_ _1061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6181_ _2111_ _2130_ _2136_ _2137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_112_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5132_ _0869_ _0874_ _0985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5063_ _0885_ _0896_ _0909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_38_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4014_ _3072_ _3174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4481__A2 _3309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5965_ _1897_ _3251_ _1900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5430__A1 _0080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5430__B2 _1311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4916_ _0745_ _0746_ _0747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_40_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5896_ _1821_ _1824_ _1825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5168__B _1023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4847_ _0663_ _0667_ _0671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4778_ _1048_ _0596_ _0602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5733__A2 _1644_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6781__I1 _2628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3729_ _2332_ _2495_ _2889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6517_ _3103_ _3185_ _2501_ _2502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6448_ _2424_ _2427_ _2428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5497__A1 _1370_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6379_ _2345_ _2352_ _2353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5631__B _1533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4472__A2 _0285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5016__A4 _2660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6858__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3432__B1 _0993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3983__A1 _3134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6772__I1 _3262_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5724__A2 _1635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3735__A1 _2893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5488__A1 _0829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4936__I _0655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4999__B1 _0837_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5660__A1 _0963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5660__B2 _1564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5750_ _1601_ _1602_ _1665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_15_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4701_ _0520_ _0524_ _0525_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5681_ _0948_ _0395_ _1589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4632_ _0449_ _0450_ _0456_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5715__A2 _0969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6763__I1 _3169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4563_ _0313_ _0387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3514_ B\[1\]\[1\] _1927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6302_ _2131_ _1811_ _2134_ _2269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4494_ _0313_ _0318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5479__A1 _1362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6233_ _2192_ _2193_ _2194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3445_ _1147_ _1158_ _1169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6164_ _1486_ _2118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4846__I _0669_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5115_ _0955_ _0956_ _0966_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6095_ _1923_ _1271_ _2043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3750__I _2849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5046_ _0621_ _0886_ _0890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_84_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4454__A2 _0277_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3662__B1 _1938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5403__A1 _3399_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5948_ _0542_ _0577_ _1880_ _1881_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3965__A1 _3115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5879_ _1584_ _1805_ _1806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_4_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6301__I _0696_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4390__A1 _0197_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4142__A1 _2945_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5890__A1 _1199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5642__A1 _1248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5945__A2 _1817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6370__A2 _2002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3835__I _2950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4381__A1 _0136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3723__A4 _1993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4133__A1 _3222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4684__A2 _0451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4666__I _0476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4436__A2 _0237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6681__I0 _2661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6851_ _0034_ net11 net1 B\[0\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5802_ _1721_ _1722_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_62_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3994_ _3147_ _3153_ _3154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6782_ _2734_ _0048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3947__A1 _3039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5733_ _1643_ _1644_ _1646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_50_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5664_ _1556_ _1559_ _1569_ _1570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_136_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4615_ _0421_ _0437_ _0438_ _0439_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5595_ _1441_ _1493_ _1494_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_50_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4546_ _0367_ _0368_ _0370_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4477_ _0246_ _0300_ _0301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6216_ _1954_ _1958_ _2174_ _2175_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3428_ _0872_ _0982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6147_ _1274_ _2099_ _2100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6078_ _2012_ _2023_ _2024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_73_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5029_ _2984_ _0870_ _0871_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5388__B1 _0585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5927__A2 _1858_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3705__A4 _2863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4115__A1 _3274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6187__B _2142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5615__A1 _1498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5918__A2 _0075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6040__A1 _1935_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3929__A1 _3078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6591__A2 _2563_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4400_ _0221_ _0222_ _0223_ _0224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5380_ _1245_ _1256_ _1258_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4331_ _0153_ _0154_ _0155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4106__A1 _3260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4262_ _3398_ _0084_ _0086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6097__B _2044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6001_ _3239_ _3284_ _1939_ _1940_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4657__A2 _3174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4396__I _3399_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4193_ _3305_ _3353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4409__A2 B\[1\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5606__A1 _1504_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6834_ _0017_ net11 net1 A\[2\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_62_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5909__A2 _1834_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6765_ _2637_ _3098_ _2719_ _2722_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5385__A3 _1262_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3977_ _3127_ _3136_ _3137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5716_ _1607_ _1626_ _1627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_137_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6696_ net10 _2673_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5647_ _1545_ _1550_ _1551_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3475__I A\[3\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4345__A1 _0107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4345__B2 _0168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5578_ _1421_ _1425_ _1475_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4896__A2 _0634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4529_ _3095_ _3383_ _0353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6098__A1 _1980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5845__A1 _0476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6270__A1 _2232_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6454__C _2421_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4820__A2 _2985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6573__A2 _2558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4584__A1 _0351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5086__B _0931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4336__A1 _3392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4887__A2 _0689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6696__I net10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4639__A2 _0408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput9 input_val[6] net9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3900_ _2596_ _2773_ _3060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4880_ _0706_ _2092_ _0708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6013__A1 _2970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3831_ _2982_ _2986_ _2987_ _2990_ _2991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_20_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6550_ _2268_ _2527_ _2534_ _1270_ net27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3762_ _0883_ _2922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5501_ _1350_ _1390_ _1391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6481_ _2456_ _2457_ _2464_ _2465_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3693_ _2799_ _2835_ _2852_ _2853_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5432_ _0164_ _0684_ _1315_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4878__A2 _2882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5363_ _2893_ _1239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3550__A2 _2310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4314_ _3345_ _1081_ _0138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5294_ _1160_ _1162_ _1163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_59_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4245_ _3379_ _0069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4176_ _3332_ _3335_ _3336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_83_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6252__A1 _1896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6004__A1 _3268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6817_ _0000_ net11 net1 A\[0\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6748_ _2663_ _0998_ _2706_ _2710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6307__A2 _0670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6679_ _2659_ _0009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4869__A2 _0687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3933__I _3006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3541__A2 _1960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6491__A1 _2401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4764__I B\[2\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5046__A2 _0886_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4557__A1 _0345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3532__A2 _2004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5809__A1 _1630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4088__A3 _3246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4030_ _3176_ _3177_ _3190_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5285__A2 _1150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5037__A2 _0876_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5981_ _1879_ _1917_ _1918_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_64_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3599__A2 _1169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4932_ _0586_ _0883_ _0765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4863_ B\[0\]\[2\] _0689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6602_ _3296_ _2581_ _2588_ _2101_ _2589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_21_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4548__A1 _0087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3814_ _2964_ _2973_ _2974_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4794_ B\[0\]\[4\] _0618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6533_ _2268_ _2511_ _2518_ _2400_ net25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3745_ _2839_ _2902_ _2905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6464_ _2442_ _2445_ _2446_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3676_ _2799_ _2835_ _2836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_133_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5415_ B\[0\]\[2\] _1296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6395_ _2173_ _2175_ _2371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5346_ _0775_ _0776_ _0831_ _0841_ _1220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_102_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5277_ _1139_ _1143_ _1144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5276__A2 _1141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4228_ _3095_ _3383_ _3387_ _1982_ _3388_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_29_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4159_ _3306_ _3316_ _3318_ _3319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_46_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4539__A1 _0331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5200__A2 _1046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4711__A1 _1785_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4494__I _0313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3838__I _2994_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput12 sel_in[0] net12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4950__A1 _2157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3530_ B\[1\]\[0\] _2102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3753__A2 _2900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3461_ A\[3\]\[6\] _1345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5200_ _1047_ _1046_ _1054_ _1060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_112_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6180_ _2132_ _2134_ _2136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_124_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5131_ _0871_ _0873_ _0984_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6455__A1 _2044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5062_ _0904_ _0906_ _0908_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_42_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4013_ _3168_ _3172_ _3173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4769__A1 _0587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5964_ _1897_ _0317_ _1898_ _1564_ _1899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5430__A2 _1310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4915_ _2515_ _0689_ _0746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3441__A1 _1037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3748__I _2907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5895_ _1556_ _1822_ _1823_ _1824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4846_ _0669_ _0670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5194__A1 _0876_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5963__I _3251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4777_ _0600_ _0883_ _0601_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4941__A1 _2790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3744__A2 _1840_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6516_ _3186_ _2453_ _2501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3728_ _2828_ _2831_ _2887_ _2888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6447_ _2346_ _2425_ _2426_ _2427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3659_ _2718_ _2746_ _2819_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6378_ _2346_ _2351_ _2352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_115_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5329_ _1200_ _3225_ _0816_ _1201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_103_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4472__A3 _0295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3680__A1 _2779_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3432__A1 _0971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3432__B2 _1015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3983__A2 _3135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3735__A2 _2894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4932__A1 _0586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4489__I _3297_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5488__A2 _0128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6437__A1 _2415_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4448__B1 _0069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4999__A1 _0836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4999__B2 _1367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5660__A2 _0133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4700_ _0521_ _0381_ _0522_ _0523_ _0515_ _0518_ _0524_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai33_1
XTAP_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5680_ _0946_ _0255_ _1588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5176__A1 _1030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4631_ _0449_ _0450_ _0455_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_129_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4562_ _0306_ _0384_ _0385_ _0386_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_6301_ _0696_ _2268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3513_ _1257_ _1268_ _1916_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4493_ _2948_ _0317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6232_ _1906_ _1914_ _2193_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3444_ B\[1\]\[3\] _1158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4687__B1 _0506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6163_ _2115_ _2117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5114_ _0962_ _0964_ _0965_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6094_ _1188_ _2039_ _2040_ _2041_ _2042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5100__A1 _0948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5045_ _0888_ _3008_ _0889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3662__B2 _2821_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5403__A2 _0618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5947_ _0544_ _0576_ _1880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3965__A2 _3124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5878_ _1586_ _1661_ _1804_ _1805_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_139_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6789__I _2731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4829_ _1367_ _0651_ _0652_ _2787_ _0653_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_21_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4914__A1 A\[2\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4102__I _2343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4142__A2 _3301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3941__I _3045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5890__A2 _1817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6825__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5642__A2 _0357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3405__A1 _0707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6699__I net13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4905__A1 _0733_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3708__A2 _0916_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4381__A2 _1004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5108__I _0837_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4133__A2 _3287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6681__I1 _0191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3644__A1 _2764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6850_ _0033_ net11 net1 B\[0\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_39_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5801_ _1717_ _1720_ _1721_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5397__A1 _3334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6781_ _1772_ _2628_ _2733_ _2734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3993_ _3148_ _3151_ _3152_ _3153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_50_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3947__A2 _3106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5732_ _1643_ _1644_ _1645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_31_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5149__A1 _1002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5663_ _1560_ _1568_ _1569_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4614_ _0424_ _0427_ _0438_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5594_ _1489_ _1492_ _1493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4545_ _0367_ _0368_ _0369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_132_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4476_ _0248_ _0299_ _0300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6558__B _2044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4857__I _0681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6215_ _1956_ _2174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3427_ _0960_ _0971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6848__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5872__A2 _1798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6146_ _2094_ _2098_ _2099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6077_ _2021_ _2022_ _2023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_39_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5028_ B\[2\]\[4\] _0870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input10_I input_val[7] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5688__I _0958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5388__A1 _3296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5388__B2 _1265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4060__A1 _2980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4899__B1 _2430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6468__B _2449_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5863__A2 _1788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5379__A1 _0857_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3846__I _1389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4354__A2 _0177_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4330_ _3274_ _2809_ _0152_ _0114_ _0154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_114_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5303__A1 _1123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4106__A2 _1235_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3581__I B\[1\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4261_ _3398_ _0084_ _0085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6000_ _3241_ _3283_ _1939_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I execute vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4192_ _3351_ _1015_ _3352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5606__A2 _1505_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6833_ _0016_ net11 net1 A\[2\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__5909__A3 _1838_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6764_ _2721_ _0041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4042__A1 _3139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3976_ _3131_ _3134_ _3135_ _3136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5715_ _0325_ _0969_ _1626_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4593__A2 _0416_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6695_ _2672_ _0014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5646_ _1546_ _1548_ _1549_ _1550_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__4345__A2 _1971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5577_ _1432_ _1445_ _1473_ _1474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5542__B2 _1287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4896__A3 _0636_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4528_ _0350_ _3032_ _3034_ _0351_ _0352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4587__I _0152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6098__A2 _1983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4459_ _2930_ _0282_ _0283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5845__A2 _1140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3856__A1 _3005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6129_ _2078_ _2079_ _2080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3608__A1 _2761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4584__A2 _0407_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5533__A1 _1421_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4336__A2 _2644_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6089__A2 _2035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3830_ _2985_ _2988_ _2922_ _2989_ _2990_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4024__A1 _3182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3761_ B\[3\]\[7\] _2921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5500_ _1293_ _1324_ _1390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6480_ _2462_ _2464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3692_ _2802_ _2834_ _2852_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5431_ _1308_ _1309_ _1313_ _1302_ _1314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_65_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4327__A2 _0148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5524__A1 _1293_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5362_ _0853_ _0860_ _1237_ _1238_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4313_ _0136_ _1004_ _0137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5293_ _1044_ _1161_ _1162_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_87_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4244_ _0064_ _0066_ _0067_ _0068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_99_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4175_ _3334_ _1389_ _3335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6816_ _2756_ _0063_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4015__A1 _3025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6747_ _2709_ _0034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3959_ _3110_ _3111_ _3119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3486__I B\[3\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6678_ _2658_ _0473_ _2656_ _2659_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5629_ _1432_ _1445_ _1531_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5515__A1 _3346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4318__A2 _0126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6491__A2 _2404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4254__A1 _2037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4006__A1 _3155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5754__A1 _3297_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4088__A4 _3247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5980_ _1881_ _1915_ _1917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_80_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4931_ _0726_ _0761_ _0763_ _0764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5993__A1 _3220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4862_ _0687_ _3271_ _0688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6601_ _1981_ _2583_ _2584_ _2587_ _2225_ _2588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_20_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3813_ _2883_ _2972_ _2973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4548__A2 _0118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4793_ _0614_ _0616_ _0617_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_119_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6532_ _2418_ _2513_ _2517_ _2518_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3744_ _1774_ _1840_ _1752_ _2904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6463_ _2371_ _2443_ _2444_ _2445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3675_ _2802_ _2834_ _2835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5414_ _0686_ _0069_ _1295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6394_ _2367_ _2369_ _2370_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_127_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5345_ _0843_ _0863_ _1218_ _1219_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5276_ _1073_ _1141_ _1142_ _1128_ _1143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_87_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4227_ _3380_ _3387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4484__A1 _0307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4158_ _3317_ _0927_ _3318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6225__A2 _1980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4089_ _2966_ _2971_ _3249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4236__A1 _3389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4814__B _0632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5200__A3 _1054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4711__A2 _0420_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4775__I B\[2\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4778__A2 _0596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput13 sel_in[1] net13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4950__A2 B\[0\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3460_ _1312_ _1323_ _1334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5130_ _0968_ _0978_ _0981_ _0983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5258__A3 _1102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5061_ _0904_ _0906_ _0902_ _0907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_84_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4466__A1 _3333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4012_ _3107_ _3170_ _3171_ _3158_ _3172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_111_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6207__A2 _1946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5963_ _3251_ _1898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5966__A1 _0290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4914_ A\[2\]\[7\] _0681_ _0745_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5894_ _1559_ _1569_ _1823_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3441__A2 _1103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4845_ _0668_ _0669_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4776_ _0599_ _0600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5194__A2 _1049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6391__A1 _2361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6515_ _2264_ _2500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3727_ _2824_ _2827_ _2887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4941__A2 _0649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6446_ _2345_ _2352_ _2426_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3658_ _2804_ _2817_ _2818_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_106_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4154__B1 _3313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6377_ _2120_ _2348_ _2350_ _2351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3589_ _2146_ _2704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5328_ _1199_ _1200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5249__A3 _1112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5259_ _1080_ _1089_ _1060_ _1124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_29_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5957__A1 _0564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3432__A2 _0982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5709__A1 _0668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6757__I0 _2673_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3735__A3 _2684_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4932__A2 _0883_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3499__A2 _1741_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6437__A2 _2300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4448__A1 _2766_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4448__B2 _1290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4999__A2 _2949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6748__I0 _2663_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4630_ _0453_ _0454_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5176__A2 _1031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4561_ _3368_ _3174_ _0385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6300_ _2103_ _2144_ _2187_ _2265_ _2266_ net21 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_3512_ _1883_ _1894_ _1905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6125__A1 _1834_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4492_ _0315_ _0316_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6231_ _1884_ _1904_ _2192_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3443_ A\[2\]\[2\] _1147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6162_ _2114_ _2115_ _2116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5113_ _0963_ _2998_ _1818_ _0959_ _0964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6093_ _0945_ _2034_ _2032_ _2041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4439__A1 _0226_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5044_ _0848_ _0888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6061__B1 _2003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5946_ _0537_ _0540_ _1878_ _1879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5877_ _1714_ _1801_ _1802_ _1803_ _1804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__6840__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4828_ _0594_ _0652_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4759_ _0527_ _0582_ _0583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4914__A2 _0681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6116__A1 _1250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6429_ _2272_ _2285_ _2407_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4602__A1 _0359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3405__A2 _0718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6831__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5158__A2 _1012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4905__A2 _0734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5330__A2 _0815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5094__A1 _0940_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5800_ _1716_ _1718_ _1720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6780_ _2731_ _2733_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5397__A2 _0615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3992_ _3062_ _3063_ _3152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_90_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5731_ _1335_ _1348_ _1644_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_95_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6822__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5149__A2 _2004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5662_ _1561_ _1567_ _1568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4613_ _0424_ _0427_ _0437_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5593_ _1490_ _1491_ _1492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4544_ _3398_ _0084_ _3377_ _0368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_128_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3580__A1 _1224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4475_ _0259_ _0298_ _0299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6214_ _2003_ _2172_ _2173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3426_ _0949_ _0960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6145_ _2095_ _2097_ _2098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6076_ _0669_ _0979_ _2022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5085__A1 _0913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5027_ _0643_ _0718_ _0869_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4832__A1 _2790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5388__A2 _0583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5929_ _1816_ _1860_ _1861_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_55_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4899__B2 _0706_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3571__A1 _2408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4115__A3 _3244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5076__A1 _0921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6328__A1 _2140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5119__I _0969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4260_ _0068_ _0083_ _0084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_125_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4191_ _3350_ _3351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4814__A1 _0634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3617__A2 _2774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6016__B1 _1378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6832_ _0015_ net11 net1 A\[1\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_91_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6763_ _2634_ _3169_ _2719_ _2721_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3975_ _3031_ _3053_ _3135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4042__A2 _3146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5714_ _1604_ _1611_ _1625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6319__A1 _2269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6694_ _2671_ _2131_ _2666_ _2672_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5645_ _0612_ _3387_ _1549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5576_ _1418_ _1431_ _1473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4527_ _0328_ _0351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3772__I _2931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4458_ _0281_ _0282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3409_ B\[3\]\[5\] _0773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4389_ _0200_ _0212_ _0213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__3856__A2 _3015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6128_ _1835_ _1837_ _2079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6059_ _1378_ _2003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4805__A1 _2810_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3608__A2 _2764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4584__A3 _0350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5781__A2 _1640_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4024__A2 _1829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6838__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3760_ _2916_ _2919_ _2920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_13_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3691_ _2847_ _2850_ _2851_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5430_ _0080_ _1310_ _1002_ _1311_ _1313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_12_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5361_ _0846_ _0852_ _1237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4312_ A\[1\]\[7\] _0136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5292_ _1154_ _1142_ _1159_ _1161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_141_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4243_ _3382_ _1158_ _0067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4174_ _3333_ _3334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6815_ _1877_ _2649_ _2751_ _2756_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4015__A2 _3174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6143__I _1865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6746_ _2661_ _1007_ _2706_ _2709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3958_ _3110_ _3111_ _3118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3774__A1 _2930_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3889_ _3047_ _3048_ _3049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6677_ net4 _2658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5515__A2 _0829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5628_ _1470_ _1518_ _1529_ _1530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4318__A3 _0141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3526__A1 _2026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5559_ _1451_ _1453_ _1454_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_105_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5931__B _1863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6779__A1 _1267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4254__A2 _0069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5451__A1 _1328_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4006__A2 _3165_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5203__A1 _1062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5754__A2 _0830_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5506__A2 _0255_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3517__A1 _1938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5690__A1 _0963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5442__A1 A\[0\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4930_ _0730_ _0736_ _0763_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5993__A2 _3218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4861_ _0686_ _0687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6600_ _1115_ _1182_ _2585_ _2587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_61_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3812_ _2966_ _2971_ _2972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4792_ _1378_ _0615_ _0616_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3756__A1 _2858_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6531_ _1162_ _2514_ _2516_ _1925_ _2517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3743_ _2839_ _2902_ _2903_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3674_ _2818_ _2833_ _2834_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6462_ _2374_ _2385_ _2444_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3508__A1 _1136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5413_ A\[0\]\[5\] _0681_ _1294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6393_ _2361_ _2366_ _2368_ _2369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5344_ _0845_ _0862_ _1218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5275_ _0980_ _1818_ _1142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4226_ _3385_ _2894_ _3386_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4484__A2 _2939_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5681__A1 _0948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4157_ A\[1\]\[3\] _3317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6582__B _2418_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4088_ _3243_ _3245_ _3246_ _3247_ _3248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_71_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4236__A2 _3395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5433__A1 _0073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3995__A1 _3115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6729_ _2696_ _0027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4172__A1 _1312_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_35 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5672__A1 _1199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5424__A1 _1299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4791__I B\[2\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6712__S _2682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5727__A2 _1343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3738__A1 _2886_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput14 sel_in[2] net14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5127__I _3005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5060_ _0675_ _1829_ _0906_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5663__A1 _1560_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4466__A2 _0773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4011_ _3015_ _1818_ _3171_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5962_ _0287_ _1897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5966__A2 _1900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4913_ _0715_ _0742_ _0743_ _0744_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5893_ _1559_ _1569_ _1822_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_33_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5718__A2 _3390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4844_ B\[2\]\[7\] _0668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3729__A1 _2332_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4775_ B\[2\]\[3\] _0599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6421__I _1269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6514_ _2400_ _2478_ _2499_ net24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3726_ _2815_ _2885_ _2886_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6445_ _2351_ _2425_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3657_ _2808_ _2816_ _2817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_106_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4154__A1 _0971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4154__B2 _3307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3588_ _1927_ _2697_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6376_ _2117_ _2240_ _2349_ _2350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5327_ _0668_ _1199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3780__I _2939_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5258_ _1057_ _1093_ _1102_ _1123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_130_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4209_ _3368_ _3369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5189_ _0961_ _1047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5406__B2 _1285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3968__A1 _3084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5709__A2 _0342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6757__I1 _2120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4393__A1 _0072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6487__B _3296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4696__A2 _0514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5893__A1 _1559_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4448__A2 _3382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5645__A1 _0612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6070__A1 _0834_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3959__A1 _3110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6748__I1 _0998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3865__I _3024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4384__A1 A\[1\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4560_ _3297_ _2940_ _0384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3511_ _1422_ _1411_ _1894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4491_ _2948_ _0313_ _0314_ _2995_ _0315_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__6125__A2 _1838_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6230_ _1912_ _1913_ _2189_ _2191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3442_ _0806_ _1114_ _1125_ _1136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4687__A2 _0459_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5884__A1 _1811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6161_ _0824_ _2115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5112_ _0836_ _0963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6092_ _1194_ _1193_ _1264_ _2040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__5636__A1 _0080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6684__I0 _2663_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5043_ _0621_ _0886_ _0887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3647__B1 _2310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5939__A2 _0524_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6061__A1 _1595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6061__B2 _2005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5945_ _1877_ _1817_ _0541_ _1878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_80_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5876_ _1662_ _1713_ _1803_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4827_ _0596_ _0651_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4375__A1 _0151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4758_ _0581_ _0582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3709_ _2867_ _2868_ _2869_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6116__A2 _0562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4689_ _0452_ _0512_ _0459_ _0513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4127__A1 _3224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6428_ _2405_ _2406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_122_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6359_ _2188_ _2329_ _2330_ _2331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6675__I0 _2652_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6052__A1 _1251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4602__A2 _0360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6871__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4905__A3 _2814_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4118__A1 _2890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4669__A2 _0492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5618__A1 _1470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5094__A2 _0941_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6043__A1 _1219_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6594__A2 _2566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3991_ _3141_ _3149_ _3150_ _3151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5730_ _1627_ _1640_ _1641_ _1643_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5661_ _1563_ _1566_ _1567_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4357__A1 _0126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4612_ _0432_ _0435_ _0436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5592_ _1222_ _0547_ _0548_ _0613_ _1491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_129_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4543_ _0349_ _0365_ _0366_ _0367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3580__A2 _1147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4474_ _0261_ _0297_ _0298_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_116_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5857__A1 _1765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6213_ _2907_ _2172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3425_ B\[3\]\[2\] _0949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6144_ _1584_ _1864_ _2096_ _2097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5609__A1 _1375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6075_ _2019_ _2020_ _2021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5026_ _0673_ _0867_ _0868_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_54_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4832__A2 _0655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6585__A2 _2453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5928_ _1826_ _1859_ _1860_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_110_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5859_ _1766_ _1780_ _1784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6337__A2 _2172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4899__A2 _0628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4115__A4 _3271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4520__A1 _0336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5076__A2 _0922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6273__A1 _1243_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6025__A1 _2946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6576__A2 _2561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4339__A1 _0148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4304__I A\[1\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6500__A2 _2448_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4511__A1 _0326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4190_ A\[1\]\[6\] _3350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6264__A1 _2226_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4814__A2 _0636_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6016__A1 _1955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6016__B2 _1898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6831_ _0014_ net11 net1 A\[1\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__6567__A2 _2544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6811__I0 _0317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6762_ _2720_ _0040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3974_ _3117_ _3132_ _3133_ _3134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5713_ _1388_ _1391_ _1624_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6693_ net9 _2671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5527__B1 _0712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5644_ _1429_ _1539_ _1547_ _1479_ _1548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_15_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5575_ _1414_ _1447_ _1471_ _1472_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4526_ _0282_ _0350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_132_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4457_ _0065_ _0281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3408_ _0740_ _0751_ _0762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4388_ _0204_ _0211_ _0212_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4884__I _0692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3856__A3 _3011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6127_ _1562_ _1836_ _2078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5058__A2 _0901_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6058_ _1955_ _2002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4805__A2 _0628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3608__A3 _2767_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5009_ _0848_ _2452_ _0849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6802__I0 _3075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4569__A1 _0392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4584__A4 _3169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3792__A2 _2951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4741__A1 _0265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4794__I B\[0\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4980__A1 _0675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3690_ _1785_ _2849_ _2850_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5574__B _1446_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3873__I _2299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4732__A1 _0551_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5360_ _1220_ _1234_ _1236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_114_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4311_ _3316_ _0132_ _0134_ _3354_ _0135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_113_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5291_ _1155_ _1159_ _1160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6485__A1 _2323_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4242_ _2343_ _0065_ _0066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4496__B1 _3368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4173_ A\[1\]\[6\] _3333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4209__I _3368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5460__A2 _1343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3471__A1 _1444_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6814_ _2755_ _0062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5212__A2 _3106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6745_ _2708_ _0033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3957_ _3006_ _3116_ _3117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3774__A2 _2933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6676_ _2657_ _0008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3888_ _2441_ _3038_ _2059_ _3048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__4879__I _0620_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5627_ _1472_ _1517_ _1529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3783__I _1532_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3526__A2 _2048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5558_ _1381_ _1452_ _1453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4509_ _3304_ _3320_ _0333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_132_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5489_ _1375_ _1371_ _1376_ _1377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_132_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6779__A2 net12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6400__A1 _2909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5203__A2 _2923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4962__A1 _2690_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4789__I _0612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5506__A3 _0128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3517__A2 _1949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4714__A1 _0285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5690__A2 _0313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5442__A2 _0627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3453__A1 _1235_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5993__A3 _3287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4860_ _0684_ _0686_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3811_ _2968_ _2970_ _2971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4791_ B\[2\]\[0\] _0615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6530_ _0388_ _0489_ _0492_ _2516_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__4953__A1 _0731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3756__A2 _2871_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3742_ _2851_ _2901_ _2902_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_9_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6461_ _2374_ _2385_ _2443_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3673_ _2820_ _2832_ _2833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_134_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5412_ _1277_ _1292_ _1293_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6392_ _0584_ _2368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5343_ _1209_ _1216_ _1217_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4181__A2 _1598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5274_ _3102_ _1140_ _1141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4225_ _3323_ _3385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5681__A2 _0395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4156_ A\[1\]\[5\] _1510_ _3316_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4087_ _3044_ _3247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5433__A2 _1296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3995__A2 _3124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4989_ _0825_ _0788_ _0792_ _0826_ _0827_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_6728_ _2663_ _3225_ _2692_ _2696_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4944__A1 _0774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6659_ _1437_ _2642_ _2638_ _2643_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4172__A2 _3328_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6449__A1 _2342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6828__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5672__A2 _0530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3683__A1 B\[3\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6492__C _2264_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5424__A2 _1303_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3688__I _0905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput15 sel_out[0] net15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4312__I A\[1\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6239__I _3245_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5143__I _0625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4010_ _3102_ _3169_ _3170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_96_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6612__A1 _0514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5961_ _1893_ _1895_ _1896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4912_ _2732_ _2821_ _0716_ _0682_ _0743_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_34_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3977__A2 _3136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5892_ _1563_ _1820_ _1821_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4843_ _0665_ _0666_ _0667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6702__I _2678_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3729__A2 _2495_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4774_ _0597_ _0993_ _0598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6513_ _2147_ _2485_ _2490_ _2491_ _2498_ _2499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3725_ _2878_ _2884_ _2885_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_20_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6444_ _2239_ _2241_ _2424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_134_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3656_ _2811_ _2815_ _2816_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5351__A1 _0855_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4154__A2 _3309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6375_ _2347_ _2160_ _2349_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3587_ A\[2\]\[6\] _2690_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5326_ _0673_ _0867_ _1197_ _1198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3901__A2 _3060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5257_ _1115_ _1121_ _1122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4208_ _3367_ _3368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3665__A1 A\[2\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5188_ _1041_ _1045_ _1046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4139_ A\[1\]\[2\] _3299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5406__A2 _1281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6813__S _2751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3968__A2 _3085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4393__A2 B\[1\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5590__B2 _1428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5893__A2 _1569_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6059__I _1378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5645__A2 _3387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3408__A1 _0740_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3959__A2 _3111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5581__A1 _0623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4384__A2 _0817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3510_ _1213_ _1279_ _1883_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4490_ _0307_ _0314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3441_ _1037_ _1103_ _1125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5884__A2 _0530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6160_ _1482_ _2114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3895__A1 _3031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5111_ _0873_ _0961_ _0962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6091_ _1194_ _1264_ _2039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5042_ _1180_ _0618_ _0886_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6684__I1 _0530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3647__A1 _2651_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3647__B2 _2806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6061__A2 _2002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5944_ _2909_ _1877_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4072__A1 _2907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5875_ _1659_ _1660_ _1802_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4826_ _1345_ _0649_ _0650_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4757_ _0529_ _0580_ _0581_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5572__A1 _0669_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3708_ _1345_ _0916_ _2868_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4688_ _0508_ _0509_ _0512_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_119_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4127__A2 _3286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6427_ _2275_ _2401_ _2404_ _2405_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_3639_ _2779_ _2795_ _2798_ _2799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_108_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6358_ _2219_ _2220_ _2218_ _2330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_143_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3886__A1 _3043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3886__B2 _3045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5309_ _1115_ _1178_ _1179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6289_ _2252_ _2254_ _2255_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6675__I1 _0491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3810__A1 _2969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4905__A4 _2810_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5315__A1 _1116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3629__B2 _2788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4054__A1 _3211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3990_ _3144_ _3145_ _3150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_62_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5660_ _0963_ _0133_ _0958_ _1564_ _1566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_128_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4611_ _0433_ _0434_ _0435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4357__A2 _0141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5591_ _0613_ _1222_ _0354_ _0357_ _1490_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_129_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4542_ _0363_ _0364_ _0366_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6839__D _0022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4473_ _0278_ _0296_ _0297_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6212_ _2156_ _2170_ _2171_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3424_ _0905_ _0927_ _0938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6143_ _1865_ _2096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6074_ _2014_ _2018_ _2020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5025_ _0810_ _0866_ _0867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_100_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6034__A2 _3285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5927_ _1828_ _1858_ _1859_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5858_ _1761_ _1782_ _1783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_16_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5545__A1 _1282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4809_ B\[0\]\[7\] _0633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5545__B2 _1319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5789_ _1647_ _1652_ _1707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_135_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3571__A3 _2535_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3859__A1 _0729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4284__A1 _0107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6025__A2 _3253_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4036__A1 _3155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5536__A1 _1311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5839__A2 _1761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4511__A2 _3015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6264__A2 _2227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6016__A2 _0317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4990__I _0599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6830_ _0013_ net11 net1 A\[1\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_36_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6811__I1 _2645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6761_ _2628_ _0407_ _2719_ _2720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3973_ _3120_ _3123_ _3133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5712_ _1618_ _1621_ _1622_ _1623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6692_ _2670_ _0013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5643_ _0561_ _0997_ _1278_ _1311_ _1547_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5527__B2 _0168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5574_ _1415_ _1325_ _1446_ _1471_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4525_ _0331_ _0348_ _0349_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4750__A2 _0573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4456_ _0204_ _0211_ _0279_ _0280_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3407_ B\[3\]\[4\] _0751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4387_ _0207_ _0210_ _0211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_58_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6126_ _1830_ _2075_ _2076_ _2077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6057_ _1999_ _2000_ _2001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6861__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5008_ B\[0\]\[5\] _0848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4018__A1 _3176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6802__I1 _2634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5766__A1 _0694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4569__A2 _0971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4405__I _0164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4741__A2 _0564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4257__A1 _0080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6731__S _2698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4980__A2 _3225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5146__I _0999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4310_ _3351_ _3307_ _2988_ _0133_ _0134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5290_ _1069_ _1157_ _1159_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4241_ _3325_ _0065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4496__A1 _0317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4496__B2 _0319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4172_ _1312_ _3328_ _3332_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5996__A1 _2981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3471__A2 _0817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6813_ _1898_ _2647_ _2751_ _2755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6796__I0 _1811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4225__I _3323_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6744_ _2658_ _1140_ _2706_ _2708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3956_ _2943_ _3116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4420__A1 _3371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6675_ _2652_ _0491_ _2656_ _2657_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3887_ _3038_ _3041_ _3042_ _3046_ _3047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__4971__A2 _0807_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5626_ _1464_ _1467_ _1527_ _1528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5920__A1 _1848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5557_ _1379_ _1383_ _1452_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4508_ _0326_ _3093_ _0331_ _0332_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5488_ _0829_ _0128_ _1376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4439_ _0226_ _0236_ _0262_ _0263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6109_ _1897_ _2058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5987__A1 _1923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6787__I0 _0830_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4962__A2 _0620_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5506__A4 _0870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4714__A2 _0295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6726__S _2692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5690__A3 _0314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3453__A2 _1246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4650__A1 _3181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3810_ _2969_ _2813_ _2267_ _2660_ _2970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_82_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4790_ _0613_ _1323_ _0614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3741_ _2853_ _2900_ _2901_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3884__I _2201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4953__A2 _2026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6460_ _2377_ _2437_ _2440_ _2442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_3672_ _2828_ _2831_ _2832_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_12_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5411_ _1286_ _1291_ _1292_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_63_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5902__A1 _1546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6391_ _2361_ _2366_ _2367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_127_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5342_ _1211_ _1215_ _1216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_142_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5273_ _1064_ _1140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_88_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4469__A1 _0291_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4224_ _3045_ _3383_ _3384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4155_ _3306_ _3310_ _3312_ _3314_ _3315_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3692__A2 _2834_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4086_ _3108_ _3246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6870__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5197__A2 _1054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4988_ _0787_ _0791_ _0826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6727_ _2695_ _0026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3939_ _3008_ _3098_ _3099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6146__A1 _2094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6658_ net7 _2642_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5609_ _1375_ _1508_ _1405_ _1406_ _1509_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6589_ _2571_ _2574_ _2575_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5121__A2 _0972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4880__A1 _0706_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3435__A2 _0850_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3986__A3 _3145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6861__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput16 sel_out[1] net16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4699__A1 _0345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4871__A1 _0689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3879__I _2113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5960_ _0273_ _0572_ _1895_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4623__A1 _0439_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4911_ _2892_ _0716_ _0682_ _2690_ _0742_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5891_ _1561_ _1567_ _1820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6852__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6376__A1 _2117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4842_ _0644_ _0647_ _0666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4773_ _0596_ _0597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4503__I A\[0\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6512_ _2492_ _2497_ _2225_ _2498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3724_ _2880_ _2881_ _2883_ _2884_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3655_ _2812_ _2813_ _2814_ _2288_ _2815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6443_ _2337_ _2355_ _2423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6374_ _2347_ _1992_ _2348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3586_ A\[2\]\[6\] _1927_ _2684_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5325_ _0810_ _0866_ _1197_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5256_ _1116_ _1119_ _1120_ _1121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_87_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4207_ _3301_ _3367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5187_ _1040_ _1044_ _1045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_130_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4862__A1 _0687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3665__A2 _1927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4138_ _2942_ _3297_ _3298_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6165__I _0562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6603__A2 _2578_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4069_ _2927_ _2976_ _3229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4614__A1 _0424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6843__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4917__A2 _0747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5342__A2 _1215_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4853__A1 _0642_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3408__A2 _0751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4605__A1 _0419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6834__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5030__A1 _0833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5581__A2 _0070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3592__A1 _2146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3440_ _1037_ _1103_ _1114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6530__A1 _0388_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5154__I _0712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5110_ _2994_ _0959_ _0961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6090_ _2027_ _2030_ _2038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5041_ _0875_ _0882_ _0884_ _0885_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3647__A2 _2660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6597__A1 _3206_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5943_ _1869_ _1870_ _1871_ _1875_ _1876_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6825__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4072__A2 _3116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6713__I _2686_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5874_ _1747_ _1799_ _1800_ _1801_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_61_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4825_ B\[2\]\[2\] _0649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5021__A1 _0845_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4233__I _3392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6818__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4756_ _0532_ _0579_ _0580_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5572__A2 _0191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3707_ A\[3\]\[7\] _0949_ _2867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4687_ _0452_ _0459_ _0506_ _0507_ _0510_ _0511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_6426_ _2276_ _2284_ _2403_ _2404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3638_ _1653_ _2796_ _2797_ _2798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5324__A2 _1195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6521__A1 _0492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3569_ _2515_ _2525_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6357_ _2219_ _2220_ _2218_ _2329_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5308_ _1174_ _1175_ _1178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6288_ _2001_ _2008_ _2253_ _2254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5239_ _1097_ _1100_ _1101_ _1102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_124_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4835__A1 _0654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_78 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6588__A1 _2572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4063__A2 _2978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3810__A2 _2813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5012__A1 _0846_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5563__A2 _1458_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5702__I _0326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3629__A2 _1059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6291__A3 _2257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6579__A1 _0506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4054__A2 _3213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5251__A1 _0873_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4610_ _0341_ _0319_ _0399_ _0434_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5590_ _1320_ _1478_ _1487_ _1428_ _1489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4541_ _0363_ _0364_ _0365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_144_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4472_ _0280_ _0285_ _0295_ _0296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_144_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6211_ _2164_ _2169_ _2170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3423_ _0916_ _0927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5857__A3 _1780_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3868__A2 _2774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6142_ _1586_ _1661_ _1804_ _1866_ _2095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_98_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6073_ _2014_ _2018_ _2019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_97_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4817__A1 _0631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5024_ _0819_ _0865_ _0866_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_39_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5490__A1 _0643_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5926_ _1839_ _1857_ _1858_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5793__A2 _1602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5857_ _1765_ _1766_ _1780_ _1759_ _1749_ _1782_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_55_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4808_ _2760_ B\[2\]\[0\] _0632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5545__A2 _1427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5788_ _1678_ _1704_ _1705_ _1706_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_4739_ _0562_ _3262_ _0563_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6409_ _2371_ _2374_ _2385_ _2386_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_116_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4808__A1 _2760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4284__A2 _1971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4036__A2 _3165_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4511__A3 _0331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5472__A1 _0651_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6760_ _2717_ _2719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5775__A2 _1628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3972_ _3120_ _3123_ _3132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3786__A1 _2945_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5711_ _1614_ _1617_ _1622_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6691_ _2669_ _1612_ _2666_ _2670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5642_ _1248_ _0357_ _1546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5527__A2 _1310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5573_ _1468_ _1469_ _1470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4524_ _0325_ _3007_ _0348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4455_ _0207_ _0210_ _0279_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3406_ A\[3\]\[2\] _0740_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4386_ _0208_ _0209_ _0210_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_59_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3710__A1 _2866_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6125_ _1834_ _1838_ _2076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6056_ _0857_ _1255_ _2000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5007_ _2525_ _0618_ _0847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5215__A1 _0918_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5766__A2 _0114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5909_ _1830_ _1834_ _1838_ _1839_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_50_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3701__A1 _2843_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5454__A1 _3323_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4257__A2 _2113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3768__A1 _2866_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4240_ _3399_ _2310_ _0064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4496__A2 _0318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4171_ _3329_ _3330_ _3331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5445__A1 _1281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6812_ _2754_ _0061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6796__I1 _2649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6743_ _2707_ _0032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3955_ _3094_ _3113_ _3114_ _3115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6721__I _2691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6674_ _2655_ _2656_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3886_ _3043_ _3040_ _3044_ _3045_ _3046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5625_ _1526_ _0191_ _1468_ _1527_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4184__A1 _3307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5556_ _1369_ _1386_ _1450_ _1451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4507_ _0330_ _0331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5487_ _3333_ _0769_ _1375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4438_ _0228_ _0235_ _0262_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4369_ _0188_ _0192_ _0193_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_115_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6108_ _1832_ _2055_ _2056_ _2057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5436__A1 _0848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6039_ _1923_ _0674_ _1981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5987__A2 _1271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3998__A1 _3097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_21 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6787__I1 _2640_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4175__A1 _3334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4151__I _3299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3922__A1 _3081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5690__A4 _0959_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5427__A1 _0102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4650__A2 _0189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6742__S _2706_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4938__B1 _0770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3740_ _2873_ _2899_ _2900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3671_ _2805_ _2829_ _2830_ _2831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_118_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6851__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5410_ _1287_ _1288_ _1289_ _1291_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_6390_ _2038_ _2042_ _2262_ _2364_ _2366_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_127_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5902__A2 _1549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5341_ _0823_ _1212_ _1214_ _1215_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5272_ _1067_ _1128_ _1130_ _1139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_142_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5666__A1 _1502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4223_ _3382_ _3383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4154_ _0971_ _3309_ _3313_ _3307_ _3314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4085_ _3244_ _3245_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4641__A2 _0416_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4987_ _0824_ _2933_ _0825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6726_ _2661_ _2910_ _2692_ _2695_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3938_ _2048_ _3098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6657_ _2641_ _0003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3869_ _3003_ _3014_ _3029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5608_ _0286_ _0878_ _1508_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6588_ _2572_ _0585_ _2573_ _2574_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5539_ _1418_ _1431_ _1432_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5657__A1 _0836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5409__A1 _0731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4880__A2 _2092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6874__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6737__S _2698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4320__A1 _0101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4871__A2 _2495_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4623__A2 _0440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4910_ _0709_ _0720_ _0739_ _0741_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5890_ _1199_ _1817_ _1819_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3831__B1 _2987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4841_ _0589_ _0664_ _0665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4772_ B\[2\]\[1\] _0596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6511_ _2421_ _2493_ _2496_ _2431_ _2497_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3723_ _1290_ _2766_ _2882_ _1993_ _2883_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6442_ _2340_ _2353_ _2422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3654_ A\[2\]\[1\] _2814_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6373_ _1239_ _2347_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6220__B _2178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3585_ _2627_ _2636_ _2668_ _2676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_138_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5324_ _0945_ _1195_ _1196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5255_ _1028_ _1029_ _1120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6300__A2 _2144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4206_ _3364_ _3365_ _3366_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5186_ _2998_ _1043_ _1044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4862__A2 _3271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4137_ A\[1\]\[0\] _3297_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4068_ _3227_ _3228_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5811__A1 _1731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4614__A2 _0427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4378__A1 A\[1\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6709_ _2683_ _0018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6678__I0 _2658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4853__A2 _0660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4605__A2 _0428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5030__A2 _1576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3592__A2 _2484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6040__B _1981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4541__A1 _0363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5040_ _0880_ _0881_ _0884_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6046__A1 _1236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5942_ _1873_ _1874_ _1875_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5873_ _1797_ _1798_ _1800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_33_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4824_ _0644_ _0647_ _0648_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5021__A2 _0862_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4755_ _0534_ _0578_ _0579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3706_ _2864_ _2792_ _2865_ _2866_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4686_ _0508_ _0509_ _0510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_135_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6425_ _2278_ _2402_ _2403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3637_ _1488_ _1554_ _2797_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6521__A2 _2226_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4532__A1 _0281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6356_ _1921_ _2222_ _2328_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3568_ A\[2\]\[6\] _2515_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5307_ _1173_ _1176_ _1177_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6287_ _2006_ _2253_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3499_ _1697_ _1741_ _1763_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5238_ _0996_ _1018_ _1101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_57_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4835__A2 _0658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6176__I _1564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5169_ _0930_ _0931_ _1025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6037__A1 _1975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6588__A2 _0585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4599__A1 _0414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3574__A2 _2565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6512__A2 _2497_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6276__A1 _1223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4826__A2 _0649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3503__I _1796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5003__A2 _0827_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4540_ _3378_ _3396_ _0364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_128_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4471_ _0288_ _0294_ _0295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6210_ _1957_ _2167_ _2169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3422_ B\[3\]\[3\] _0916_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6141_ _2089_ _2093_ _2094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_124_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6072_ _2016_ _2017_ _2018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5023_ _0821_ _0864_ _0865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6019__A1 _1956_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5490__A2 _0307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5925_ _1842_ _1856_ _1857_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_34_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5856_ _1765_ _1766_ _1780_ _1781_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_22_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4807_ _0619_ _0621_ _0624_ _0630_ _0631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5787_ _1702_ _1703_ _1705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4738_ _0561_ _0562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4669_ _0489_ _0492_ _0493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4505__A1 _0328_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6408_ _2379_ _2384_ _2385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_122_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6339_ _2306_ _2307_ _2308_ _2309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4808__A2 B\[2\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3492__A1 _1433_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5769__B1 _0546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3795__A2 _2936_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4992__A1 _2938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4744__A1 _0073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4511__A4 _0333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5472__A2 _3317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3483__A1 _1565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5224__A2 _1001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4027__A3 _3186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3971_ _3129_ _3130_ _3131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5710_ _1619_ _1621_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6690_ net8 _2669_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5641_ _0824_ _1223_ _0547_ _0548_ _1545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_86_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5572_ _0669_ _0191_ _1469_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4523_ _0324_ _0334_ _0347_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4454_ _0263_ _0277_ _0278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_102_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5160__A1 _0975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3405_ _0707_ _0718_ _0729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4385_ A\[1\]\[6\] _0916_ _0209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6124_ _1834_ _1838_ _2075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_98_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3710__A2 _2869_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6055_ _1252_ _1254_ _1999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5006_ _0745_ _0746_ _0799_ _0801_ _0846_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_38_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4974__A1 _0760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5908_ _1835_ _1837_ _1838_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_14_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5839_ _1760_ _1761_ _1762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3701__A2 _2860_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4149__I _3308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5454__A2 _0690_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5206__A2 _0800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4965__A1 _3260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3768__A2 _2869_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4717__A1 _0537_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5142__A1 _0975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4170_ _3324_ _3326_ _3330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_67_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6642__A1 net2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5445__A2 _1326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6811_ _0317_ _2645_ _2751_ _2754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_63_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6742_ _2652_ _1731_ _2706_ _2707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3954_ _3104_ _3112_ _3114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6673_ _2630_ _2654_ _2655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3885_ _2113_ _3045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5624_ _1200_ _1526_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5381__A1 _1238_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4184__A2 _3313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5555_ _1370_ _1385_ _1450_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4506_ _3326_ _0329_ _0330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3931__A2 _3078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5486_ _1371_ _1372_ _1373_ _1364_ _1374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_105_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4437_ _0214_ _0238_ _0260_ _0261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5353__I _0586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4368_ _2921_ _0191_ _0192_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3695__A1 _2789_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6107_ _1852_ _1853_ _2056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4299_ _3349_ _3355_ _0123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6633__A1 _1195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5436__A2 _0220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6038_ _1935_ _1979_ _1980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_100_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3998__A2 _3103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4947__A1 _0760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4432__I _0255_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5372__A1 _1247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4175__A2 _1389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5372__B2 _1248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5124__A1 _3005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5675__A2 _1581_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6624__A1 _2225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5427__A2 _0692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3438__A1 _1070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3989__A2 _3145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4938__B2 _1356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3670_ _1224_ _1993_ _2830_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4166__A2 _2310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5340_ _0827_ _0842_ _1214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_115_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3913__A2 _3072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5115__A1 _0955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5271_ _1131_ _1132_ _1127_ _1138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_99_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4222_ A\[0\]\[3\] _3382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4153_ _3305_ _3313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6615__A1 _3211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5418__A2 _1295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4084_ _2879_ _3244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4517__I _0318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3421__I _0740_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6732__I _2699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4929__A1 _0730_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4986_ _0613_ _0824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3937_ _2932_ _3096_ _3097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6725_ _2694_ _0025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5348__I _1221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3601__A1 _2760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6656_ _0548_ _2640_ _2638_ _2641_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3868_ _1872_ _2774_ _3028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5607_ _1503_ _1506_ _1507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6587_ _1173_ _1176_ _2573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3799_ _2525_ _1191_ _2959_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5538_ _1426_ _1430_ _1431_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5469_ _1353_ _1354_ _1355_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_105_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5657__A2 _3334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5409__A2 _0327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6082__A2 _1262_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output25_I net25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5345__A1 _0843_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3659__A1 _2718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4320__A2 _0117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3831__A1 _2982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4840_ _0590_ _0828_ _0664_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4771_ _1048_ _0594_ _0595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6510_ _2424_ _2427_ _2494_ _1923_ _2496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3722_ A\[2\]\[2\] _2882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5336__A1 _1199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6441_ _2356_ _2360_ _2421_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3653_ _2765_ _2813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6372_ _1243_ _1996_ _2243_ _2244_ _2249_ _2346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_3584_ _2651_ _2660_ _2668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5323_ _1188_ _1193_ _1194_ _1195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5254_ _1108_ _1117_ _1118_ _1119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4956__B _0790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4205_ _3359_ _3363_ _3365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5185_ _1042_ _1043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4136_ _3295_ _3296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4067_ _2916_ _2919_ _3226_ _3227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4075__A1 _2936_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5811__A2 _0351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3822__A1 _2786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4378__A2 B\[3\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4969_ _0783_ _0804_ _0805_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6708_ _2661_ _3246_ _2682_ _2683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6639_ _2101_ _2622_ _2625_ _2626_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_137_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3889__A1 _3047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6678__I1 _0473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4853__A3 _0611_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4066__A1 _2908_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6841__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5015__B1 _2092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6358__A3 _2218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5566__A1 _1394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5318__A1 _0907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5869__A2 _1715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6530__A3 _0492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6748__S _2706_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4541__A2 _0364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4829__B1 _0652_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5941_ _0244_ _0301_ _0529_ _0580_ _1874_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_80_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3804__A1 _2958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5872_ _1797_ _1798_ _1799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_55_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4823_ _0645_ _0646_ _0647_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_21_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5557__A1 _1379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4754_ _0542_ _0577_ _0578_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3705_ _2760_ _1356_ _1510_ _2863_ _2865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_105_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4685_ _0501_ _0500_ _0509_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4530__I _3385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6424_ _2283_ _2402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3636_ _1488_ _1554_ _2796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6521__A3 _2503_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6355_ _0520_ _2324_ _2325_ _2326_ _2327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3567_ _2484_ _2495_ _2505_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4532__A2 _3098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5306_ _1174_ _1175_ _1176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_89_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6286_ _1200_ _2003_ _2252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3498_ _1697_ _1741_ _1752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_103_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5237_ _1082_ _1098_ _1099_ _1100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6457__I _2383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6864__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4296__A1 _0087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5493__B1 _0255_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5168_ _0994_ _1022_ _1023_ _1024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6037__A2 _1978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4119_ _3276_ _3278_ _3279_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_17_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5099_ _0597_ _0948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4599__A2 _0415_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3810__A4 _2660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4771__A2 _0594_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5720__A1 _0065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5539__A1 _1418_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5003__A3 _0842_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4470_ _0289_ _0293_ _0294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_128_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3421_ _0740_ _0905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6140_ _2090_ _2091_ _2093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6071_ _1230_ _1232_ _2017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5181__I _0878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5475__B1 _1360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5022_ _0843_ _0863_ _0864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_85_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5778__A1 _1691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5924_ _1847_ _1855_ _1856_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_62_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5855_ _1768_ _1775_ _1778_ _1779_ _1780_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_139_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4806_ _0626_ _0629_ _0630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5786_ _1702_ _1703_ _1704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4737_ _0168_ _0561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4668_ _0490_ _0491_ _0407_ _0472_ _0492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3619_ _1422_ _2771_ _2778_ _2779_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4505__A2 _3032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6407_ _2380_ _2383_ _2384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4599_ _0414_ _0415_ _0423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6338_ _2172_ _2306_ _2308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6269_ _2012_ _2023_ _2233_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5769__A1 _0281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5769__B2 _1068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4441__A1 _0079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3795__A3 _2954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4992__A2 _0830_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4744__A2 _2969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5941__B2 _0580_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3704__B1 _2863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3483__A2 _1576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6761__S _2719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3970_ _3000_ _3001_ _3130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_51_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6560__I _1267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5640_ _1537_ _1542_ _1544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6185__A1 _2139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5571_ _1464_ _1467_ _1468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_79_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4522_ _3374_ _0119_ _0346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4453_ _0269_ _0276_ _0277_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3404_ A\[3\]\[0\] _0718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5160__A2 _1001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4384_ A\[1\]\[7\] _0817_ _0208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6123_ _2054_ _2073_ _2074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6054_ _1990_ _1997_ _1998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_112_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5999__A1 _3234_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5005_ _0793_ _0803_ _0844_ _0845_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4671__A1 _0388_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4423__A1 _0195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5907_ _1562_ _1836_ _1837_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_22_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5838_ _1725_ _1742_ _1743_ _1761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_139_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5769_ _0281_ _1064_ _0546_ _1068_ _1685_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5151__A2 _3246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6645__I _2631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4165__I A\[0\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4414__A1 _0216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4965__A2 _0800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5914__A1 _0888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6714__I0 _2669_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3940__A3 _3097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6642__A2 net12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4653__A1 _0476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6810_ _2752_ _0060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6741_ _2705_ _2706_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_51_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3953_ _3104_ _3112_ _3113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6504__B _2488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4803__I B\[0\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6672_ net2 _2653_ _2654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3884_ _2201_ _3044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4708__A2 _0253_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5905__A1 _1229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5623_ _1522_ _1524_ _1525_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3419__I _0872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5554_ _1392_ _1448_ _1449_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_144_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4505_ _0328_ _3032_ _0329_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6705__I0 _2658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5485_ _1363_ _1358_ _1373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_144_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4436_ _0216_ _0237_ _0260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4367_ _0190_ _0191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3695__A2 _2793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6106_ _1854_ _2055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4298_ _3349_ _3355_ _0122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6633__A2 _0585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6037_ _1975_ _1978_ _1979_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_67_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6873__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_78 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5124__A2 _0970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6624__A2 _2610_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3438__A2 _1081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6864__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4938__A2 _0769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5060__A1 _0675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5270_ _1124_ _1135_ _1137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_99_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5115__A2 _0956_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4221_ _3037_ _3380_ _3381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3677__A2 _2836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4152_ _3311_ _0927_ _3312_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6615__A2 _3213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4083_ _2930_ _3243_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6855__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4929__A2 _0736_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4985_ _0768_ _0778_ _0822_ _0823_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5051__A1 _0893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4533__I _0149_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6724_ _2658_ _1829_ _2692_ _2694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3936_ _3095_ _3096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3601__A2 _1389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6655_ net6 _2640_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3867_ _3023_ _3026_ _3021_ _3027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5606_ _1504_ _1505_ _1506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4689__B _0459_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6586_ _1173_ _1176_ _2572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3798_ _2825_ _2826_ _2891_ _2895_ _2958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_118_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5537_ _1427_ _1428_ _1429_ _1430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_133_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6303__A1 _2111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5468_ _0590_ A\[1\]\[1\] _1354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4419_ _0180_ _0241_ _0243_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5399_ _0627_ _1278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4865__A1 _0690_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3668__A2 _2827_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6846__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4093__A2 _2950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5290__A1 _1069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3840__A2 _2999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5042__A1 _1180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output18_I net18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3659__A2 _2746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6837__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5033__A1 _0651_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4770_ B\[2\]\[2\] _0594_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3595__A1 _2684_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3721_ _2812_ _2806_ _2881_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6440_ _2414_ _2416_ _2418_ _2420_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6533__A1 _2268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3652_ _2762_ _2812_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5336__A2 _1208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3583_ _1949_ _2660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6371_ _2342_ _2344_ _2345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5184__I _0651_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5322_ _0868_ _0944_ _1194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_142_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5253_ _1111_ _1112_ _1118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_102_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4204_ _3359_ _3363_ _3364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5184_ _0651_ _1042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4135_ _3288_ _3295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4066_ _2908_ _3225_ _2920_ _3226_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_113_38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6828__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4075__A2 _2954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5272__A1 _1067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6743__I _2707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5811__A3 _0350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3822__A2 _0982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4968_ _0793_ _0803_ _0804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_71_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6707_ _2678_ _2682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_138_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3919_ _2996_ _3079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4899_ _2967_ _0628_ _2430_ _0706_ _0728_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6524__A1 _2500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6638_ _2623_ _2624_ _2625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6569_ _3199_ _2147_ _2553_ _2554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3889__A2 _3048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4838__A1 _0642_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6819__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4066__A2 _3225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5263__A1 _1067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5015__A1 _0734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5015__B2 _0733_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4173__I A\[1\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3577__A1 _2473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6602__B _2588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4901__I _0633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4829__A1 _1367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5940_ _0529_ _0580_ _1873_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3804__A2 _2963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5871_ _1712_ _1706_ _1710_ _1798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__4083__I _2930_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4822_ _0590_ _1070_ _0646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4753_ _0544_ _0576_ _0577_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6512__B _2225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3704_ _2760_ _1510_ _2863_ _1499_ _2864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_105_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4684_ _0444_ _0451_ _0508_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6423_ _2116_ _2121_ _2401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3635_ _2783_ _2794_ _2795_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3427__I _0960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6354_ _1873_ _1874_ _2326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_127_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3566_ A\[2\]\[4\] _2495_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5305_ _1124_ _1135_ _1123_ _1175_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_103_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6285_ _2237_ _2250_ _2251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3497_ _1719_ _1730_ _1741_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5236_ _1085_ _1088_ _1099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4296__A2 _0118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5493__B2 _0837_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5167_ _1020_ _1021_ _1023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_97_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4118_ _2890_ _3261_ _3277_ _2960_ _3278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5098_ _0946_ _0982_ _0947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5245__A1 _1100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4048__A2 _3152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4049_ _3148_ _3208_ _3209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5796__A2 _1703_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5720__A2 _0690_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6648__I net4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5484__A1 _0597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4168__I A\[0\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5787__A2 _1703_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3420_ _0861_ _0883_ _0894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6070_ _0834_ _1231_ _2016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_48_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5475__A1 _1358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input9_I input_val[6] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5021_ _0845_ _0862_ _0863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_79_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5778__A2 _1694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5923_ _1832_ _1854_ _1855_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_94_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5854_ _1768_ _1775_ _1779_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4805_ _2810_ _0628_ _0629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5785_ _1625_ _1645_ _1703_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4736_ _0229_ _3033_ _0560_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4667_ _0341_ _0491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6406_ _2200_ _2381_ _2382_ _2383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6831__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3618_ _2759_ _2770_ _2778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4598_ _0414_ _0415_ _0422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6337_ _2058_ _2172_ _2307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3549_ _2299_ _2310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6268_ _1989_ _2011_ _2232_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5466__A1 _0586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5219_ _1063_ _1078_ _1079_ _1080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6199_ _1943_ _1950_ _2155_ _2156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5769__A2 _1064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4441__A2 _2299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6718__A1 _2649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4744__A3 _2766_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3952__A1 _3009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3704__A1 _2760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3704__B2 _1499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5209__A1 _1068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3530__I B\[1\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6185__A2 _2140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6854__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5570_ _1396_ _1465_ _1467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3943__A1 _3101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4521_ _0340_ _0343_ _0344_ _0345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4452_ _0223_ _0275_ _0276_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5696__A1 _0327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3403_ B\[3\]\[6\] _0707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4383_ _0205_ _0138_ _0206_ _0207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6122_ _2064_ _2072_ _2073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6053_ _1243_ _1996_ _1997_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_85_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5004_ _0796_ _0802_ _0844_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4120__A1 _2970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4423__A2 _0239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5906_ _0287_ _0959_ _1836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5837_ _1749_ _1759_ _1760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4187__A1 _3346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5768_ _3328_ _1007_ _1684_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3934__A1 _3093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4719_ _0263_ _0277_ _0543_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5699_ _0325_ _0969_ _1607_ _1608_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_136_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5439__A1 _1318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4414__A2 _0237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6661__I net8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6877__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4965__A3 _0711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6167__A2 _2120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5914__A2 _1482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6714__I1 _2160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3525__I _2037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4653__A2 _3169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5850__A1 _1771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6772__S _2724_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6740_ _2629_ _2703_ _2705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3952_ _3009_ _3110_ _3111_ _3112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_44_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6671_ net12 _2653_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3883_ _2070_ _3043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4169__A1 _3262_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4091__I _0707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5622_ _1523_ _1519_ _1524_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5905__A2 _0326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3916__A1 _2994_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5553_ _1414_ _1447_ _1448_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_129_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4504_ _0327_ _0328_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5484_ _0597_ _0128_ _1372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6705__I1 _2933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5669__A1 _1503_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4435_ _0254_ _0258_ _0259_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4341__A1 _0164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4366_ _0189_ _0190_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6105_ _1839_ _1857_ _2053_ _2054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4297_ _3374_ _0119_ _0120_ _0121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6036_ _3228_ _1976_ _1977_ _1978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6633__A3 _2619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_35 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6869_ _0052_ net11 net1 B\[2\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__5097__I _0770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4580__A1 _0328_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5124__A3 _0975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4332__A1 _0151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4883__A2 _0681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6085__A1 _1198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4399__A1 _2969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5060__A2 _1829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5899__A1 _1553_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6767__S _2719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4220_ _3379_ _3380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4151_ _3299_ _3311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6076__A1 _0669_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4082_ _2867_ _2868_ _2941_ _2953_ _3242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_110_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4086__I _3108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4984_ _0774_ _0777_ _0822_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6723_ _2693_ _0024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3935_ _3037_ _3095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6654_ _2639_ _0002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3866_ _2921_ _3025_ _3026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5605_ _3346_ _0870_ _1505_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6585_ _2569_ _2453_ _2570_ _2571_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3797_ _2886_ _2897_ _2956_ _2957_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5536_ _1311_ _0997_ _1429_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5467_ A\[1\]\[2\] _0588_ _1353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4418_ _0180_ _0241_ _0242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5398_ _1275_ _1276_ _1277_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4865__A2 _2806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4349_ _0163_ _0172_ _0173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_86_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4617__A2 _0439_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6019_ _1956_ _1958_ _1959_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5042__A2 _0618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4305__A1 _0128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5033__A2 _0982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3720_ _2879_ _2288_ _2880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4792__A1 _1378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3651_ _2809_ _2354_ _2810_ _1301_ _2811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6533__A2 _2511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6370_ _0670_ _2002_ _2341_ _2344_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3582_ _2644_ _2651_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5321_ _1189_ _1034_ _1190_ _1192_ _1184_ _1186_ _1193_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai33_1
XFILLER_142_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5252_ _1111_ _1112_ _1117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_88_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4847__A2 _0667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4203_ _3361_ _3362_ _3363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5183_ _0950_ _1038_ _1040_ _1041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_111_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6049__A1 _1250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4134_ _0696_ _3293_ _3294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4065_ _2923_ _3225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5811__A4 _1140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4967_ _0796_ _0802_ _0803_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_52_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3586__A2 _1927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6706_ _2681_ _0017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4783__A1 _0600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3918_ _3074_ _3077_ _3078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4898_ _0627_ _1949_ _0727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6637_ _3221_ _3291_ _2624_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3849_ _3008_ _2961_ _3009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6568_ _3193_ _3198_ _2553_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5519_ _1374_ _1377_ _1410_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6499_ _2449_ _2447_ _2482_ _2483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6288__A1 _2001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4838__A2 _0660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3577__A2 _2545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4774__A1 _0597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6602__C _2101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4829__A2 _0651_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6451__A1 _2422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5870_ _1762_ _1747_ _1764_ _1794_ _1795_ _1797_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_34_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4821_ _0588_ _1532_ _0645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4752_ _0557_ _0575_ _0576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4765__A1 _1070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3703_ _0949_ _2863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4683_ _0500_ _0503_ _0507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6422_ _2268_ _2301_ _2399_ _2400_ net22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_135_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3634_ _2789_ _2793_ _2794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_128_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6353_ _0302_ _0524_ _0581_ _2325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__5190__A1 _0652_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3565_ B\[1\]\[2\] _2484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5304_ _1106_ _1113_ _1174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_89_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3740__A2 _2899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6284_ _2244_ _2249_ _2250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3496_ _1587_ _1642_ _1730_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5235_ _1085_ _1088_ _1098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5493__A2 _0392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5166_ _1020_ _1021_ _1022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_112_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6754__I _2714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4117_ _2959_ _2962_ _3277_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_99_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5097_ _0770_ _0946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5245__A2 _1101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4048_ _3151_ _3152_ _3208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5999_ _3234_ _3237_ _1936_ _1937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4508__A1 _0326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5484__A2 _0128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5989__B _1925_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6664__I net9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4995__A1 _0833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4747__A1 _0233_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3528__I A\[2\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6672__A1 net2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5020_ _0853_ _0860_ _0862_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5899__B _1827_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5922_ _1852_ _1853_ _1854_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_34_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5853_ _1667_ _1776_ _1777_ _1778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__6523__B _2101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4804_ _0627_ _0628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5784_ _1680_ _1700_ _1701_ _1702_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4735_ _0269_ _0276_ _0558_ _0559_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3410__A1 _0773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3961__A2 _3036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4666_ _0476_ _0490_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6405_ _2240_ _2198_ _2349_ _2382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_135_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6749__I _2710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3617_ _1872_ _2774_ _2776_ _2777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4597_ _3007_ _0420_ _0421_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6336_ _2206_ _2207_ _1900_ _2306_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3548_ B\[1\]\[4\] _2299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6267_ _2021_ _2022_ _2019_ _2231_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3479_ _1081_ _1532_ _1543_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4269__A3 A\[0\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5218_ _1071_ _1077_ _1079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6198_ _1951_ _1961_ _2155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3477__A1 _1499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5149_ _1002_ _2004_ _1003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5218__A2 _1077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4729__A1 _0286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3401__A1 net16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4744__A4 _3380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3952__A2 _3110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3704__A2 _1510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3468__A1 _1334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5209__A2 _3035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6406__A1 _2200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4968__A1 _0793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3640__A1 _2616_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5393__A1 _3295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5932__A3 _1863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4520_ _0336_ _0339_ _0344_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3943__A2 _3102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4451_ _0271_ _0274_ _0275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_117_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3402_ _0685_ _0696_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5696__A2 _0972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4382_ _0136_ _3333_ _1004_ _0960_ _0206_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6121_ _2065_ _2071_ _2072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_124_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5448__A2 _1276_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6052_ _1251_ _1995_ _1996_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_86_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5003_ _0823_ _0827_ _0842_ _0843_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_26_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5620__A2 _1458_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5905_ _1229_ _0326_ _1835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3631__A1 _2790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5836_ _1758_ _1759_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4187__A2 _2786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5767_ _1068_ _0411_ _1683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4718_ _0535_ _0541_ _0542_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3934__A2 _2923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5698_ _1606_ _1607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4649_ _3369_ _0473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6319_ _2269_ _2286_ _2287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_131_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6636__A1 _3220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3870__A1 _3004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5611__A2 _1511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4462__I A\[1\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3925__A2 _3080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4886__B1 _0713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4350__A2 _0173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3861__A1 _3017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6821__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3951_ _2015_ _3105_ _3042_ _3111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_63_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3613__A1 _2616_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6670_ net3 _2652_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3882_ _2931_ _2894_ _3042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5621_ _1459_ _1460_ _1449_ _1523_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4169__A2 _3328_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5366__A1 _1241_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5552_ _1416_ _1446_ _1447_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3916__A2 _3075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4503_ A\[0\]\[0\] _0327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6299__I _1269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5483_ _3345_ _0770_ _1371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4434_ _1785_ _0257_ _0258_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4341__A2 _1938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4365_ _3311_ _0189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6104_ _2052_ _1856_ _2053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4296_ _0087_ _0118_ _0120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6035_ _3231_ _3285_ _1977_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3451__I _1224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3852__A1 _3005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6762__I _2720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3604__A1 _2762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6868_ _0051_ net11 net1 B\[2\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5357__A1 _0834_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5819_ _1737_ _1738_ _1740_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6799_ _2744_ _2745_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_109_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4580__A2 _3098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3626__I _0817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6609__A1 _2593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4457__I _0065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6085__A2 _1263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4096__A1 _3250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6844__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5832__A2 _1734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6388__A3 _2258_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4399__A2 _2813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5288__I _1062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4020__A1 _3167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3536__I B\[1\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5520__A1 _1374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4874__A3 _0700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4150_ _3307_ _3309_ _3310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6076__A2 _0979_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4367__I _0190_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4081_ _2955_ _2975_ _3240_ _3241_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5036__B1 _2943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4983_ _0781_ _0805_ _0820_ _0821_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6722_ _2652_ _3025_ _2692_ _2693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3934_ _3093_ _2923_ _3094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5339__A1 _0827_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6653_ _0547_ _2637_ _2638_ _2639_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3865_ _3024_ _3025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5604_ _1380_ _3313_ _1504_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4011__A1 _3015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6584_ _3201_ _3204_ _2570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3796_ _2888_ _2896_ _2956_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5535_ _0848_ _0088_ _1428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4562__A2 _0384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5466_ _0586_ A\[1\]\[0\] _1352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4417_ _0193_ _0240_ _0241_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_105_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4314__A2 _1081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5511__A1 _1375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5397_ _3334_ _0615_ _1276_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6867__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4348_ _0167_ _0171_ _0172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_141_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4279_ _0102_ _2398_ _0103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4078__A1 _3234_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6018_ _2946_ _1957_ _1958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4617__A3 _0440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5814__A2 _1734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5578__A1 _1421_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4250__A1 _0073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4002__A1 _3104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4553__A2 _0371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6667__I net10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4305__A2 _0751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4792__A2 _0615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6518__B1 _0472_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3650_ _1147_ _2810_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3581_ B\[1\]\[3\] _2644_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4544__A2 _0084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5320_ _0991_ _1032_ _1035_ _1033_ _1192_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_142_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5251_ _0873_ _1047_ _1107_ _1116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_47_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4202_ _3339_ _3342_ _3362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5182_ _1807_ _1039_ _1040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6049__A2 _3263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4133_ _3222_ _3287_ _3292_ _3293_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4064_ _2912_ _2979_ _3223_ _3224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4966_ _0799_ _0801_ _0802_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6705_ _2658_ _2933_ _2679_ _2681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3917_ _3073_ _3076_ _3077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4783__A2 _0993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4897_ _0634_ _0725_ _0726_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6636_ _3220_ _3215_ _3218_ _2623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3848_ _1246_ _3008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6688__S _2666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6567_ _2538_ _2544_ _2552_ net28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3779_ _1081_ _2939_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5518_ _1399_ _1408_ _1409_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6498_ _2446_ _2481_ _2482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5391__I _1269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5449_ _1277_ _1332_ _1333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5799__A1 _0318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6460__A2 _2437_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output23_I net23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5971__A1 _0551_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4774__A2 _0993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5723__A1 _1295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6203__A2 _3245_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4820_ _0643_ _2985_ _0644_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4751_ _0559_ _0574_ _0575_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_1690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4765__A2 _0588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3702_ _2859_ _2861_ _2862_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4682_ _0499_ _0505_ _0506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6421_ _1269_ _2400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3633_ _2784_ _2791_ _2792_ _2793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__5714__A1 _1604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6352_ _0303_ _0582_ _2324_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3564_ _2408_ _2441_ _2212_ _2463_ _2473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_108_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5190__A2 _2984_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5303_ _1123_ _1152_ _1172_ _1173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6283_ _2007_ _2248_ _2249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_89_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3495_ _1708_ _0762_ _1719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5234_ _1095_ _1096_ _1097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5165_ _0913_ _0928_ _1021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_124_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4116_ _3273_ _3275_ _3276_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5096_ _0868_ _0944_ _0945_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_84_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4047_ _3147_ _3206_ _3207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6442__A2 _2353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5998_ _1877_ _1208_ _3238_ _1936_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5953__A1 _0561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4949_ _0738_ _0754_ _0782_ _0783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4290__I _3399_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6619_ _0514_ _0519_ _2605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4508__A2 _3093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6753__I0 _2669_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3731__A3 _2890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3495__A2 _0762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4444__A1 _0265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6680__I net5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6613__C _2264_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4747__A2 _0560_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6744__I0 _2658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5172__A2 _1025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5921_ _1480_ _1843_ _1541_ _1538_ _1853_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_34_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5852_ _1720_ _1777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4803_ B\[0\]\[4\] _0627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5783_ _1698_ _1699_ _1701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4734_ _0264_ _0268_ _0558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6735__I0 _2671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4665_ _0479_ _0488_ _0489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_134_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6404_ _2347_ _1945_ _2381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3616_ _2586_ _2775_ _2773_ _2776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5163__A2 _1017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4596_ _3353_ _0420_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6335_ _2303_ _2304_ _2305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3547_ A\[2\]\[2\] _2288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6112__A1 _1562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3478_ A\[3\]\[4\] _1532_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6266_ _2031_ _2035_ _2229_ _2230_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4269__A4 A\[0\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5217_ _1071_ _1077_ _1078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6197_ _2152_ _2153_ _2154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3477__A2 _1510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5148_ _0693_ _1002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6415__A2 _2180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5079_ _0680_ _0702_ _0926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4426__A1 _0200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6179__A1 _2060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4729__A2 _0751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6726__I0 _2661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3952__A3 _3111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3468__A2 _1400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4665__A1 _0479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4968__A2 _0803_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3640__A2 _2757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5917__A1 _1247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3539__I _2190_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5917__B2 _1222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5393__A2 _1271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4450_ _0272_ _0273_ _0274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3401_ net16 _0674_ _0685_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4381_ _0136_ _1004_ _0960_ _3350_ _0205_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_125_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6120_ _1845_ _2069_ _2071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6051_ _1244_ _1994_ _1995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4656__A1 _0472_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5002_ _0831_ _0841_ _0842_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_78_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4408__A1 _2332_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4959__A2 _0747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5081__A1 _0925_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5904_ _1545_ _1550_ _1833_ _1834_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3631__A2 _0850_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5835_ _1751_ _1756_ _1757_ _1758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6581__A1 _2566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5766_ _0694_ _0114_ _1682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4717_ _0537_ _0540_ _0541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6708__I0 _2661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5697_ _1326_ _1605_ _1606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4648_ _3182_ _0472_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4579_ _3015_ _0257_ _0403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6318_ _2272_ _2285_ _2286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6249_ _2196_ _2210_ _2211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3912__I _2988_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6876__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3870__A2 _3006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5072__A1 _0800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5375__A2 _1251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3925__A3 _2987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4886__A1 _0710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6867__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5063__A1 _0885_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3950_ _3105_ _3107_ _3109_ _3099_ _3110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_44_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3613__A2 _2757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3881_ _3039_ _3040_ _3041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5620_ _1457_ _1458_ _1454_ _1522_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5551_ _1432_ _1445_ _1446_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_77_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4502_ _0325_ _0326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6315__A1 _2120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5482_ _1327_ _1330_ _1332_ _1277_ _1370_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_144_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4326__B1 _3033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4433_ _0256_ _0257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4364_ _0183_ _0187_ _0188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6529__B _2043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6618__A2 _0518_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6103_ _1842_ _2052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4828__I _0594_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3732__I A\[2\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4295_ _0087_ _0118_ _0119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6034_ _3231_ _3285_ _1976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6858__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3852__A2 _3007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5659__I _3334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4563__I _0313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3604__A2 _2763_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6867_ _0050_ net11 net1 B\[2\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5818_ _1737_ _1738_ _1739_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6798_ _1267_ _2653_ _2730_ _2744_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_136_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5749_ _1651_ _1654_ _1663_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3540__A1 _2048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6609__A2 _2453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4738__I _0561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6849__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5293__A1 _1044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5832__A3 _1727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5045__A1 _0888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4399__A3 _3323_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4020__A2 _3179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5520__A2 _1377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4648__I _3182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3552__I _2332_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4080_ _2957_ _2974_ _3240_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5036__A1 _0878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5036__B2 _0597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4982_ _0783_ _0804_ _0820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6721_ _2691_ _2692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_108_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3933_ _3006_ _3093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6652_ _2631_ _2638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5339__A2 _0842_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3864_ _2998_ _3024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6536__A1 _1163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5603_ _1228_ _0256_ _1503_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6583_ _3201_ _3204_ _2569_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3795_ _2929_ _2936_ _2954_ _2955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_121_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5534_ _0112_ _0628_ _1427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5465_ _1293_ _1324_ _1351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4416_ _0195_ _0239_ _0240_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5511__A2 _1371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5396_ _1247_ _3328_ _1275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3522__A1 _1982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4347_ _0106_ _0169_ _0170_ _0171_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4278_ A\[0\]\[6\] _0102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5275__A1 _0980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6773__I _2727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6017_ _1955_ _1898_ _1957_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5389__I net2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5027__A1 _0643_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4250__A2 _2697_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4002__A2 _3112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5750__A2 _1602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5852__I _1720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5502__A2 _1350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3513__A1 _1257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4069__A2 _2976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6683__I net6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5018__A1 _0855_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6518__A1 _0490_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6518__B2 _0491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3580_ _1224_ _1147_ _2636_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5250_ _1106_ _1113_ _1115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4201_ _3300_ _3360_ _3361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6794__S _2738_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5181_ _0878_ _1039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4132_ _3222_ _3287_ _3291_ _3292_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4063_ _2914_ _2978_ _3223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5009__A1 _0848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6221__A3 _2178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4965_ _3260_ _0800_ _0711_ _0801_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6704_ _2680_ _0016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6509__A1 _2342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3916_ _2994_ _3075_ _3076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4896_ _0632_ _0634_ _0636_ _0725_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5980__A2 _1915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6635_ _0304_ _0525_ _2621_ _2622_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3847_ _3006_ _3007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3457__I _1290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6834__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6566_ _2546_ _2551_ _2552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3778_ _2937_ _2938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5732__A2 _1644_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3743__A1 _2839_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6768__I _2723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5517_ _1403_ _1407_ _1408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_133_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6497_ _2377_ _2479_ _2480_ _2481_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5448_ _1275_ _1276_ _1332_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5496__A1 _1374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4288__I _0111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5379_ _0857_ _1255_ _1256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_59_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5799__A2 _1043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5420__A1 _1296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3982__A1 _3134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5723__A2 _1629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5487__A1 _3333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6739__A1 net14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5411__A1 _1286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6857__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4750_ _0566_ _0573_ _0574_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3973__A1 _3120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3701_ _2843_ _2860_ _2861_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_144_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4681_ _0500_ _0504_ _0505_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6420_ _1273_ _2336_ _2370_ _2397_ _2399_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_31_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3632_ _1048_ _0916_ _2792_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6351_ _2317_ _2322_ _2323_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_115_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3563_ _2452_ _2419_ _2070_ _2430_ _2463_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5302_ _1167_ _1171_ _1172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_143_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6282_ _2246_ _2247_ _2248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3494_ _1620_ _0872_ _1708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5478__A1 _1363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5233_ _0965_ _0966_ _1096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_97_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4150__A1 _3307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5164_ _0996_ _1018_ _1019_ _1020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4115_ _3274_ _3269_ _3244_ _3271_ _3275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_68_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5095_ _0907_ _0942_ _0943_ _0944_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4046_ _3202_ _3203_ _3206_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5650__A1 _1509_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5402__A1 _0161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4205__A2 _3363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5997_ _3215_ _1930_ _1931_ _1934_ _1935_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XPHY_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4571__I _0392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4948_ _0741_ _0753_ _0782_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5953__A2 _1301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4879_ _0620_ _0706_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6618_ _0515_ _0518_ _2604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4508__A3 _0331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6753__I1 _1241_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3716__A1 _2387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6549_ _0498_ _2528_ _2533_ _2534_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3650__I _1147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5641__A1 _0824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6744__I1 _1140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3707__A1 A\[3\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3825__I _2984_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4132__A1 _3222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6357__B _2218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5880__A1 _1470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5920_ _1848_ _1850_ _1852_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5851_ _0341_ _1039_ _1776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4802_ _0625_ _2967_ _0626_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4199__A1 _3322_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5782_ _1698_ _1699_ _1700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5935__A2 _1867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4733_ _0545_ _0556_ _0557_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4664_ _3182_ _0473_ _0488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6735__I1 _2003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5699__A1 _0325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6403_ _3266_ _1948_ _2163_ _2164_ _2169_ _2380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_3615_ _1905_ _2576_ _2775_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4595_ _0403_ _0417_ _0418_ _0419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6334_ _2211_ _2216_ _2304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3546_ _2267_ _1158_ _2277_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6265_ _2027_ _2030_ _2229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_130_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6112__A2 _2061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3477_ _1499_ _1510_ _1521_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4123__A1 _3257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5216_ _0973_ _1075_ _1076_ _1077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_130_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6196_ _1963_ _1972_ _2153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5871__A1 _1712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5147_ _2933_ _0998_ _1000_ _3035_ _1001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3470__I A\[3\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5078_ _0914_ _0923_ _0924_ _0925_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input15_I sel_out[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4029_ _3172_ _3184_ _3186_ _3188_ _3189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_53_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3937__A1 _2932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6726__I1 _2910_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5862__A1 _1731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5614__A1 _1502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6662__I0 _2118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5090__A2 _0936_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5917__A2 _1486_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6590__A2 _2575_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3400_ net15 _0674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4380_ _0201_ _0203_ _0204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_131_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4105__A1 _3262_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6050_ _1991_ _1992_ _1994_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_86_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input7_I input_val[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5001_ _0832_ _0840_ _0841_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_100_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4656__A2 _0473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5853__A1 _1667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4408__A2 _3379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5605__A1 _3346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6653__I0 _0547_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5081__A2 _0926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5903_ _1548_ _1831_ _1832_ _1833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_34_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5834_ _1754_ _1755_ _1757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5765_ _1062_ _0420_ _1681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6581__A2 _1925_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4716_ _0280_ _0538_ _0539_ _0540_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6708__I1 _3246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5696_ _0327_ _0972_ _1605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4647_ _0464_ _0465_ _0462_ _0471_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__3465__I B\[3\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4578_ _0390_ _0400_ _0402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_116_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6317_ _2276_ _2284_ _2285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3529_ _2081_ _2092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6248_ _2205_ _2209_ _2210_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6636__A3 _3218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4647__A2 _0465_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5844__A1 _1754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6179_ _2060_ _2133_ _2134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3607__B1 _1180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5072__A2 _3108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4280__B1 _3037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6324__A2 _2292_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4886__A2 _0711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6686__I net7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6088__A1 _1195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6260__A1 _2188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4810__A2 _0633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3880_ _2810_ _3040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5550_ _1436_ _1443_ _1445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_117_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4501_ _0133_ _0325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5481_ _1357_ _1366_ _1368_ _1369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4326__A1 _2961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4432_ _0255_ _0256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4326__B2 _0149_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4363_ _0185_ _0186_ _0187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6079__A1 _1987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6102_ _1826_ _1859_ _2050_ _2051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4294_ _0099_ _0101_ _0117_ _0118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_98_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6033_ _1937_ _1974_ _1975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_113_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4844__I B\[2\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3852__A3 _3011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3604__A3 A\[2\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6866_ _0049_ net11 net1 B\[2\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6003__A1 _3257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5817_ _1691_ _1694_ _1681_ _1738_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_6797_ _2743_ _0055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5748_ _1623_ _1657_ _1662_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_135_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5679_ _1583_ _1585_ _1586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_117_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6609__A3 _2594_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3540__A2 _2201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5817__A1 _1691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6490__A1 _2401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4399__A4 _0161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4703__B _0526_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6545__A2 _3191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5753__B1 _0953_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5808__A1 _0282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5284__A2 _1151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5036__A2 _2922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4981_ _0816_ _0818_ _0819_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_51_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4795__A1 _2201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6720_ _2654_ _2677_ _2691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3932_ _3091_ _3092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6651_ net5 _2637_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3863_ _3021_ _3022_ _3023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5602_ _1500_ _1501_ _1502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6582_ _2564_ _2567_ _2418_ _2568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3794_ _2941_ _2953_ _2954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5533_ _1421_ _1425_ _1426_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5464_ _1335_ _1348_ _1349_ _1350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_105_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4415_ _0214_ _0238_ _0239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5395_ _1273_ _1274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4346_ _0107_ _0079_ _2102_ _2697_ _0170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__3522__A2 _2004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4277_ _0068_ _0083_ _0100_ _0101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6016_ _1955_ _0317_ _1378_ _1898_ _1956_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3899__B _3058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5027__A2 _0718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6224__A1 _1975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4786__A1 _0605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6849_ _0032_ net11 net1 B\[0\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_126_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4538__A1 _0359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5266__A2 _1077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4777__A1 _0600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3828__I _2786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6518__A2 _0407_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4200_ _2945_ _3317_ _3360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5180_ _0718_ _0951_ _1038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4131_ _3290_ _3291_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6454__A1 _2361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4062_ _2981_ _3221_ _3222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5009__A2 _2452_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4964_ _0690_ _0800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6703_ _2652_ _3102_ _2679_ _2680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3915_ _2989_ _3075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4895_ _0679_ _0722_ _0723_ _0724_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3440__A1 _1037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6634_ _0304_ _0525_ _1924_ _2621_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5717__B1 _1000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3846_ _1389_ _3006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5193__A1 _1049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6565_ _1793_ _1781_ _2550_ _0696_ _2551_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_3777_ _2790_ _2937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5516_ _1405_ _1406_ _1407_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3743__A2 _2902_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6496_ _2437_ _2440_ _2480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5447_ _1327_ _1330_ _1331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5496__A2 _1377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5378_ _1252_ _1254_ _1255_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_59_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4329_ _2809_ _0152_ _3385_ _3274_ _0153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_59_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5248__A2 _1022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5420__A2 _0111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3982__A2 _3135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5487__A2 _0769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5239__A2 _1100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5103__I _0946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3670__A1 _1224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3700_ _1444_ B\[3\]\[4\] _2860_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4680_ _0501_ _0503_ _0504_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3631_ _2790_ _0850_ _2791_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5175__A1 _1030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6350_ _2191_ _2319_ _2320_ _2322_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3562_ _2387_ _2452_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5301_ _1123_ _1170_ _1171_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6281_ _1251_ _1995_ _2247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3493_ _1136_ _1675_ _1686_ _1697_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5478__A2 _1358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5232_ _1094_ _1055_ _1095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3489__A1 _1587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5163_ _1016_ _1017_ _1019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4150__A2 _3309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6427__A1 _2275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4114_ _2969_ _3274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5094_ _0940_ _0941_ _0943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4045_ _3201_ _3204_ _3205_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4989__A1 _0825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6109__I _1897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5996_ _2981_ _1932_ _1933_ _1934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5402__A2 _0625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4947_ _0760_ _0780_ _0781_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_138_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3964__A2 _3120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4878_ _0622_ _2882_ _0705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6617_ _2147_ _2602_ _2500_ _2603_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3829_ _1015_ _2989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3716__A2 B\[1\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6548_ _2529_ _2530_ _2532_ _1273_ _2533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_134_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6479_ _2308_ _2458_ _2461_ _2462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_133_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6418__A1 _2391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5641__A2 _1223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5157__A1 _0688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3707__A2 _0949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4937__I _0649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4132__A2 _3287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3891__A1 _3011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6824__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3643__A1 _2761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5850_ _1771_ _1773_ _1775_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4801_ B\[0\]\[3\] _0625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5396__A1 _1247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5781_ _1627_ _1640_ _1699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_61_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4732_ _0551_ _0555_ _0556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_9_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4663_ _0471_ _0486_ _0487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3614_ _2596_ _2773_ _2774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6402_ _2377_ _2378_ _2379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5699__A2 _0969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4594_ _0409_ _0416_ _0418_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3545_ _2190_ _2267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6333_ _2196_ _2210_ _2303_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4371__A2 _0176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6264_ _2226_ _2227_ _2228_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3476_ B\[3\]\[1\] _1510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5215_ _0918_ _1072_ _1008_ _1076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__5320__A1 _0991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6195_ _1942_ _1962_ _2152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5146_ _0999_ _1000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3882__A1 _2931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5077_ _0921_ _0922_ _0924_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4028_ _3076_ _3187_ _3188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_72_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3634__A1 _2789_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5979_ _1906_ _1914_ _1915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_100_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3937__A2 _3096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6639__A1 _2101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5311__A1 _1116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6847__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5862__A2 _0476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6662__I1 _2645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5588__I _0075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4492__I _0315_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4050__B2 _3209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6640__C _1269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5550__A1 _1436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4353__A2 _0176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6368__B _2007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5000_ _0835_ _0838_ _0840_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5853__A2 _1776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5605__A2 _0870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6653__I1 _2637_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5902_ _1546_ _1549_ _1832_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_34_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5369__A1 _1240_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5833_ _1754_ _1755_ _1756_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4041__A1 _3199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5764_ _1679_ _1680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6550__C _1270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4715_ _0285_ _0295_ _0539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4592__A2 _0414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5695_ _1594_ _1603_ _1604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4646_ _0469_ _0470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_107_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5541__A1 _1288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4577_ _0390_ _0400_ _0401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6316_ _2278_ _2283_ _2284_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3528_ A\[2\]\[4\] _2081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6097__A2 _2042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3459_ _1246_ _1323_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6247_ _1900_ _2208_ _2209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_77_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6178_ _2057_ _2062_ _2133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5129_ _0979_ _0980_ _0975_ _0977_ _0981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_85_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3607__A1 _2766_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3607__B2 _1290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4280__A1 _0080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4280__B2 _3393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5780__A1 _1681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3791__B1 _2950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5532__A1 _1423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4271__A1 _0092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4810__A3 A\[2\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6012__A2 _3278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4023__A1 _3107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3566__I A\[2\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4500_ _0312_ _0323_ _0324_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5480_ _1362_ _1365_ _1368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4431_ _3308_ _0255_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4326__A2 _0070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5523__A1 _1307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4362_ _0127_ _0130_ _0186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6101_ _1828_ _1858_ _2050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4293_ _0110_ _0116_ _0117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6032_ _1940_ _1973_ _1974_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3837__A1 _0784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5730__B _1641_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6865_ _0048_ net11 net1 B\[2\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5816_ _1727_ _1735_ _1736_ _1737_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6796_ _1811_ _2649_ _2738_ _2743_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4565__A2 _0388_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5747_ _1659_ _1660_ _1661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5762__A1 _1599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5678_ _1520_ _1525_ _1585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5514__A1 _1401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5691__I _1599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4629_ _0316_ _0322_ _0435_ _0453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5817__A2 _1694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6490__A2 _2404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4005__A1 _3157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5087__B _0934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5753__A1 _0948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5753__B2 _3367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4308__A2 _2863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5808__A2 _1064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4980_ _0675_ _3225_ _0818_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3931_ _3079_ _3078_ _3086_ _3091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__4795__A2 _0618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5992__A1 _3220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6650_ _2635_ _0001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3862_ _3017_ _3020_ _3022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5601_ _1436_ _1443_ _1501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6581_ _2566_ _1925_ _2567_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6792__I0 _1595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3793_ _2944_ _2952_ _2953_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_121_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5532_ _1423_ _1424_ _1425_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5463_ _1346_ _1347_ _1349_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4414_ _0216_ _0237_ _0238_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5394_ _1272_ _1273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4345_ _0107_ _1971_ _2697_ _0168_ _0169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4276_ _0077_ _0082_ _0100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6015_ _2938_ _1955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6224__A2 _1978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4786__A2 _0608_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6848_ _0031_ net11 net1 A\[3\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_10_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4538__A2 _0360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5735__A1 _1350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6779_ _1267_ net12 _2730_ _2731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__6783__I0 _1043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4226__A1 _3385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5974__A1 _0552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4777__A2 _0883_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5726__A1 _1607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6774__I0 _2647_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3844__I _2949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4701__A2 _0524_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4130_ _3288_ _3289_ _3290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4061_ _3215_ _3218_ _3220_ _3221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4465__A1 _2942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4963_ _0785_ _0797_ _0798_ _0799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__5965__A1 _1897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6702_ _2678_ _2679_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3914_ _2986_ _3071_ _3073_ _3074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_71_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4894_ _0704_ _0721_ _0723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3440__A2 _1103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6633_ _1195_ _0585_ _2619_ _2620_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5717__A1 _0411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6765__I0 _2637_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5717__B2 _0328_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3845_ _3004_ _3005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6564_ _2547_ _2548_ _2549_ _2550_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3776_ _2934_ _2880_ _2885_ _2935_ _2936_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_121_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5515_ _3346_ _0829_ _1406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6495_ _2437_ _2440_ _2479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5446_ _1328_ _1329_ _1330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5377_ _0798_ _1240_ _1253_ _0849_ _1254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_87_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4328_ _3325_ _0152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4259_ _0077_ _0082_ _0083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_75_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6880__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5956__A1 _0568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6381__A1 _2337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6133__A1 _0669_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3498__A2 _1741_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4495__I _2995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5239__A3 _1101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6436__A2 _2292_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3670__A2 _1993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6215__I _1956_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3630_ A\[3\]\[7\] _2790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6372__A1 _1243_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5175__A2 _1031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3561_ _2419_ _2430_ _2441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5300_ _1137_ _1151_ _1168_ _1170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6124__A1 _1834_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6280_ _1244_ _1994_ _2246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3492_ _1433_ _1664_ _1686_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5478__A3 _1364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5231_ _1052_ _1053_ _1094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5162_ _1016_ _1017_ _1018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_123_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4113_ _1312_ _3270_ _3244_ _3272_ _3273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6427__A2 _2401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5093_ _0940_ _0941_ _0942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_112_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4044_ _3202_ _3203_ _3204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_68_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3749__I _2908_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5995_ _3224_ _3286_ _1933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_24_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3949__B1 _3108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4946_ _0764_ _0779_ _0780_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4877_ _0680_ _0702_ _0703_ _0704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6616_ _3070_ _2601_ _2602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6363__A1 _1925_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3828_ _2786_ _2988_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6547_ _1166_ _2368_ _2531_ _2532_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3759_ _2917_ _2918_ _2919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3484__I B\[3\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6115__A1 _1847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6478_ _2309_ _2314_ _2460_ _2461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5429_ _3392_ _1311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6418__A2 _2394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5204__I _1009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5641__A3 _0547_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output21_I net21 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6830__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5157__A2 _1003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4668__A1 _0490_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3891__A2 _3036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5093__A1 _0940_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3643__A2 _2764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4840__A1 _0590_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4800_ _0623_ _2931_ _0624_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5396__A2 _3328_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5780_ _1681_ _1695_ _1696_ _1698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4731_ _0552_ _0554_ _0555_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6821__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4662_ _0480_ _0485_ _0486_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6401_ _2002_ _1877_ _2375_ _2378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3613_ _2616_ _2757_ _2772_ _2773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__5699__A3 _1607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4593_ _0409_ _0416_ _0417_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_122_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6332_ _2213_ _2215_ _2302_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3544_ _1916_ _2234_ _2245_ _2256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6263_ _2188_ _1922_ _2222_ _2227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_131_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3475_ A\[3\]\[6\] _1499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4659__A1 _3182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6548__C _1273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5214_ _1072_ _1073_ _1074_ _1066_ _1075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_130_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6194_ _1969_ _1970_ _2150_ _2151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5145_ _0628_ _0999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3882__A2 _2894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5076_ _0921_ _0922_ _0923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_37_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4027_ _3183_ _3171_ _3186_ _3187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_77_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3634__A2 _2793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5978_ _1912_ _1913_ _1914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_40_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4929_ _0730_ _0736_ _0761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5139__A2 _0932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4898__A1 _0627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4103__I _2821_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6639__A2 _2622_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3942__I _3035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6879__RN net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5862__A3 _1772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5075__A1 _0710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4773__I _0596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4822__A1 _0590_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6575__A1 _1793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4050__A2 _3205_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6327__A1 _2142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5109__I _0958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3561__A1 _2419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4656__A4 _0479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4813__A1 _0632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5901_ _1546_ _1549_ _1831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5832_ _1733_ _1734_ _1727_ _1755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_62_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5763_ _1665_ _1676_ _1679_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_124_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4714_ _0285_ _0295_ _0538_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6318__A1 _2272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4592__A3 _0415_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5694_ _1601_ _1602_ _1603_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4329__B1 _3385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4645_ _0460_ _0468_ _0469_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_135_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4576_ _0391_ _0399_ _0400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_144_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6315_ _2120_ _2280_ _2282_ _2283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3527_ _1938_ _2070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3762__I _0883_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6246_ _2206_ _2207_ _2208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3458_ _1301_ _1312_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6177_ _2131_ _0670_ _2132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5128_ _0970_ _0980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5059_ _0902_ _0903_ _0904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3607__A2 A\[2\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4280__A2 _2419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4032__A2 _3191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6309__A1 _2273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3791__A1 _2948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3791__B2 _1367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5532__A2 _1424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3543__A1 _2135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4099__A2 _2973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5296__A1 _1163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5048__A1 _0614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4810__A4 _1180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5548__B _1441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5220__A1 _0970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3847__I _3006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4023__A2 _3170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5771__A2 _1682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4430_ _0250_ _0253_ _0254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6720__A1 _2654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5523__A2 _1322_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4361_ _3341_ _0184_ _0185_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3582__I _2644_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6100_ _1821_ _1824_ _2047_ _2049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4292_ _0089_ _0113_ _0115_ _0116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_98_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5287__A1 _1154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6031_ _1963_ _1972_ _1973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_112_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3837__A2 _2996_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5039__A1 _0880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4262__A2 _0084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6864_ _0047_ net11 net1 B\[1\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5815_ _1733_ _1734_ _1736_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6795_ _2742_ _0054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5211__A1 _1009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6837__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5746_ _1522_ _1524_ _1660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_136_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5677_ _1520_ _1525_ _1583_ _1584_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4628_ _0444_ _0451_ _0452_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_68_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5514__A2 _1404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4559_ _0381_ _0382_ _0383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5278__A1 _3024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6229_ _1908_ _1911_ _2189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5817__A3 _1681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6778__A1 net14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4272__B _0092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5753__A2 _0395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3764__A1 _2921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5505__A2 _3311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3616__B _2773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5269__A1 _1127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3819__A2 _2978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5441__A1 _1293_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3930_ _3089_ _3090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_45_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5992__A2 _3287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3861_ _3017_ _3020_ _3021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_32_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5600_ _1439_ _1442_ _1500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6580_ _0506_ _0507_ _0510_ _2566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3792_ _2947_ _2951_ _2952_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6792__I1 _2645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5531_ _0079_ _1296_ _1424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5462_ _1346_ _1347_ _1348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_133_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4413_ _0226_ _0236_ _0237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_132_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5393_ _3295_ _1271_ _1272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4180__A1 _0773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4344_ A\[0\]\[6\] _0168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4275_ _3336_ _0098_ _0099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_87_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6014_ _1952_ _1953_ _1954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5680__A1 _0946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6572__B _2368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5432__A1 _0164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6847_ _0030_ net11 net1 A\[3\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6778_ net14 net13 _2730_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6783__I1 _2634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3746__A1 _2904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5729_ _1638_ _1639_ _1641_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5423__A1 _1282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4226__A2 _2894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3985__A1 _3029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5726__A2 _1628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6774__I1 _2198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4021__I _3093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4060_ _2980_ _3219_ _3220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_110_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4465__A2 _3353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5414__A1 _0686_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4962_ _2690_ _0620_ _0798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5965__A2 _3251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6701_ _2629_ _2677_ _2678_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3913_ _1807_ _3072_ _3073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4893_ _0704_ _0721_ _0722_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6632_ _1194_ _1188_ _1193_ _2619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
X_3844_ _2949_ _3004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5717__A2 _0998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6765__I1 _3098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6563_ _1784_ _1792_ _2549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3775_ _2878_ _2884_ _2935_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6390__A2 _2042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5514_ _1401_ _1404_ _1405_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_118_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6494_ _2413_ _2472_ _2476_ _2477_ _2478_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_118_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5445_ _1281_ _1326_ _1329_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_105_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5376_ _0847_ _0851_ _1253_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_99_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4327_ _0067_ _0148_ _0150_ _0115_ _0151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_99_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3770__I _1312_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4258_ _0074_ _0078_ _0081_ _0082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_75_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5653__A1 _1441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4189_ _3344_ _3347_ _3348_ _3318_ _3349_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_43_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5405__A1 _0623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6381__A2 _2355_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6133__A2 _1612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4695__A2 _0518_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4776__I _0599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4447__A2 _0265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5644__B2 _1479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3958__A1 _3110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3855__I _3007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3560_ _2081_ _2430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6124__A2 _1838_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3491_ _1433_ _1664_ _1675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5230_ _1061_ _1090_ _1091_ _1093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6387__B _2258_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5161_ _0914_ _0923_ _1017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_97_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4112_ _3271_ _3272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6427__A3 _2404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5092_ _0677_ _0808_ _0941_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_84_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5635__A1 _1241_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4043_ _3196_ _3194_ _3203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5994_ _3224_ _3286_ _1932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_52_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3949__A1 _2931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3949__B2 _3045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4945_ _0768_ _0778_ _0779_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4610__A2 _0319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4876_ _0697_ _0701_ _0703_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6615_ _3211_ _3213_ _2593_ _2601_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3827_ _1796_ _0927_ _2987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6363__A2 _2334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4374__A1 _0151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6546_ _1153_ _1165_ _2531_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3758_ _2859_ _2861_ _2918_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6477_ _2311_ _2459_ _2460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3689_ _2848_ _2849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5428_ _0716_ _1310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4596__I _3353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5359_ _1227_ _1233_ _1234_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_134_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5641__A4 _0548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6051__A1 _1244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4117__A1 _2959_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5865__A1 _1718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4668__A2 _0491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3876__B1 _3034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6409__A3 _2385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3628__B1 _2786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5093__A2 _0941_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3643__A3 _2767_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4840__A2 _0828_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4730_ _0290_ _0553_ _0554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4661_ _0482_ _0484_ _0485_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6400_ _2909_ _2375_ _2377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3612_ _1422_ _2771_ _2772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6870__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4592_ _0329_ _0414_ _0415_ _0416_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_128_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6331_ _2298_ _2300_ _2301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3543_ _2135_ _2223_ _2245_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6262_ _3295_ _2225_ _2226_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3474_ _1455_ _1466_ _1092_ _1477_ _1488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_88_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5856__A1 _1765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4659__A2 _3369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5213_ _1009_ _3106_ _3040_ _1005_ _1074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6193_ _1965_ _1968_ _2150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_97_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5144_ _0997_ _0998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5608__A1 _0286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6656__I0 _0548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5075_ _0710_ _0915_ _0691_ _0922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__5084__A2 _0931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6281__A1 _1251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4026_ _3103_ _3185_ _3186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_77_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5977_ _1612_ _2908_ _1913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4928_ _0654_ _0658_ _0759_ _0760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_78 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4859_ B\[0\]\[0\] _0684_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5544__B1 _0999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4898__A2 _1949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6529_ _1044_ _1161_ _2043_ _2514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3570__A2 _1971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5847__A1 _1732_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5862__A4 _0342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5075__A2 _0915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4822__A2 _1070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4586__A1 _3043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6327__A2 _2139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4338__A1 _2343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6710__S _2682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4889__A2 _0716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3561__A2 _2430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4964__I _0690_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6263__A1 _2188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4813__A2 _0634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5900_ _1508_ _1511_ _1560_ _1568_ _1830_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_34_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6880_ _0063_ net11 net1 B\[3\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_34_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5831_ _1156_ _0190_ _1753_ _1754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_22_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5762_ _1599_ _1677_ _1678_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4713_ _0291_ _0536_ _0537_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5693_ _1592_ _1593_ _1602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6318__A2 _2285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4329__A1 _2809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4329__B2 _3274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4644_ _0462_ _0466_ _0467_ _0468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4575_ _0397_ _0398_ _0399_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6559__C _2500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3526_ _2026_ _2048_ _2059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6314_ _2117_ _2119_ _2281_ _2282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6245_ _0568_ _1889_ _2207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3457_ _1290_ _1301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5035__I _0652_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6176_ _1564_ _2131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5127_ _3005_ _0979_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5057__A2 _0901_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5058_ _0898_ _0901_ _0903_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input13_I sel_in[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4009_ _3096_ _3169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6006__A1 _3263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6557__A2 _1151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4114__I _2969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3791__A2 _2949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3543__A2 _2223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4740__A1 _0230_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6493__A1 _2300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6485__B _2468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5048__A2 _0616_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6245__A1 _0568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5220__A2 _3116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4731__A1 _0552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4360_ _1620_ A\[1\]\[4\] _0184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4291_ _1235_ _0114_ _0115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6030_ _1969_ _1970_ _1972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_112_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5287__A2 _1142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I input_val[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6236__A1 _0564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6863_ _0046_ net11 net1 B\[1\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_62_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5814_ _1733_ _1734_ _1735_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6794_ _2005_ _2647_ _2738_ _2742_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5211__A2 _3108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5745_ _1623_ _1657_ _1658_ _1659_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5676_ _1528_ _1582_ _1583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_135_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4627_ _0446_ _0449_ _0450_ _0451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__3773__I _2932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4558_ _0180_ _0241_ _3371_ _0382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_132_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3509_ _1862_ _1872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4489_ _3297_ _0313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5278__A2 _1039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6228_ _1918_ _1920_ _2188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6159_ _1845_ _2069_ _2112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6227__A1 _2147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6778__A2 net13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4109__I _2704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3948__I _2882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4961__A1 _0622_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3764__A2 _2923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4713__A1 _0291_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3860_ _3018_ _3019_ _3020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3791_ _2948_ _2949_ _2950_ _1367_ _2951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4952__A1 _0708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5530_ _0164_ _0693_ _1423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5461_ _1304_ _1305_ _1347_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3593__I A\[2\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4412_ _0228_ _0235_ _0236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__3507__A2 _1840_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5392_ _3289_ _1271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4343_ _0165_ _0166_ _0167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_141_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4274_ _0091_ _0097_ _0098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_99_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4468__B1 _2950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6013_ _2970_ _3279_ _1953_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5680__A2 _0255_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3994__A2 _3153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6846_ _0029_ net11 net1 A\[3\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6777_ _2729_ _0047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3989_ _3144_ _3145_ _3149_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5728_ _1638_ _1639_ _1640_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_108_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5659_ _3334_ _1564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6448__A1 _2424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5423__A2 _1283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3985__A2 _3057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3737__A2 _2896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5111__A1 _0873_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6827__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3673__A1 _2820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4870__B1 _0691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6611__A1 _1183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5414__A2 _0069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4961_ _0622_ _1949_ _0797_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3588__I _1927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6700_ net14 _2675_ _2677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3912_ _2988_ _3072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3976__A2 _3134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4892_ _0709_ _0720_ _0721_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_32_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6631_ _1805_ _2617_ _2618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5178__A1 _0940_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3843_ _2993_ _3002_ _3003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3728__A2 _2831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4925__A1 _0724_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6562_ _1766_ _1780_ _2548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3774_ _2930_ _2933_ _2934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5513_ _0136_ _0655_ _1404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6493_ _2300_ _2414_ _2477_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5444_ _0623_ _0327_ _1328_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5350__A1 _0824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5375_ _1249_ _1251_ _1252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4326_ _2961_ _0070_ _3033_ _0149_ _0150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3900__A2 _2773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5102__A1 _1796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4257_ _0080_ _2113_ _0081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4188_ _3306_ _3316_ _3348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_132_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6602__A1 _3296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5405__A2 _0065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6829_ _0012_ net11 net1 A\[1\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4392__A2 _0174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5644__A2 _1539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3655__A1 _2812_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3958__A2 _3111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4080__A1 _2957_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4907__A1 _0730_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5580__A1 _1311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5128__I _0970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3591__B1 _2711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3490_ _1488_ _1554_ _1653_ _1664_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_143_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5160_ _0975_ _1001_ _1013_ _1014_ _1016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_116_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3894__A1 _3051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4111_ _2081_ _3271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5091_ _0908_ _0937_ _0939_ _0940_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_97_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4042_ _3139_ _3146_ _3202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5635__A2 _1486_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5993_ _3220_ _3218_ _3287_ _1931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__4207__I _3301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3949__A2 _3043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4944_ _0774_ _0777_ _0778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_80_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4875_ _0697_ _0701_ _0702_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_60_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6614_ _2103_ _2592_ _2595_ _2600_ _2266_ net32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3826_ _2983_ _2985_ _2986_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6363__A3 _2335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6545_ _3180_ _3191_ _2145_ _2530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3757_ _2843_ _2860_ _2917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6476_ _2313_ _2459_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3688_ _0905_ _2848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5427_ _0102_ _0692_ _1309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5358_ _1230_ _1232_ _1233_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4309_ _3345_ _0133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5289_ _1156_ _3024_ _1157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3637__A1 _1488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4062__A1 _2981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3956__I _2943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5562__A1 _0668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5314__A1 _1119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4668__A3 _0407_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3876__A1 _2932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3876__B2 _3035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6708__S _2682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6665__I1 _2647_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6042__A2 _1215_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4053__A1 _3148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3800__A1 _1224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4660_ _0475_ _0483_ _0484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_119_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3611_ _2759_ _2770_ _2771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4591_ _3384_ _0410_ _0356_ _0415_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_128_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6330_ _2295_ _2297_ _2293_ _2300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3542_ _2135_ _2223_ _2234_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_116_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5305__A1 _1124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6261_ _0674_ _2225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3473_ _1059_ _0839_ _1477_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_115_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5212_ _1005_ _3106_ _1073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_88_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4659__A3 _0479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6192_ _1937_ _1974_ _2149_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5143_ _0625_ _0997_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5608__A2 _0878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6656__I1 _2640_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5074_ _0915_ _0918_ _0919_ _0920_ _0921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_56_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3619__A1 _1422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4025_ _3024_ _3181_ _3185_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4044__A1 _3202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5976_ _1908_ _1911_ _1912_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_52_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4927_ _0648_ _0659_ _0759_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4858_ _2157_ _0682_ _0683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5544__A1 _0972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3809_ B\[1\]\[6\] _2969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5544__B2 _0357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4789_ _0612_ _0613_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6528_ _3188_ _3291_ _2512_ _2513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6459_ _2380_ _2438_ _2439_ _2440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_134_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3858__A1 _0762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4807__B1 _0624_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5075__A3 _0691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4035__A1 _3167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4586__A2 _3385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4338__A2 _0161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5535__A1 _0848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4510__A2 _0333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6237__I _3243_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4274__A1 _0091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4813__A3 _0636_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5830_ _1729_ _1732_ _1753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4026__A1 _3103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5761_ _1665_ _1676_ _1677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4712_ _0289_ _0293_ _0536_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5692_ _1597_ _1600_ _1601_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5526__A1 _1318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4329__A2 _0152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4643_ _0464_ _0465_ _0467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4574_ _3310_ _0393_ _0308_ _0398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_6313_ _2279_ _2118_ _2281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3525_ _2037_ _2048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4220__I _3379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6244_ _0565_ _1888_ _2206_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3456_ B\[1\]\[6\] _1290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6175_ _2125_ _2129_ _2130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_112_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5126_ _0976_ _0977_ _0978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_111_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5057_ _0898_ _0901_ _0902_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4265__A1 _0088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4008_ _3100_ _3158_ _3160_ _3168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__5986__I net16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6006__A2 _3274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5765__A1 _1062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5959_ _0569_ _0571_ _1893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6811__S _2751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4740__A2 _1235_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6493__A2 _2414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6860__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4008__A1 _3100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6181__A1 _2111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4290_ _3399_ _0114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4247__A1 _1982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5995__A1 _3224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6862_ _0045_ net11 net1 B\[1\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_81_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5813_ _1605_ _1687_ _1688_ _1734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_62_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6793_ _2741_ _0053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5744_ _1655_ _1656_ _1658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5675_ _1530_ _1581_ _1582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6430__I _2269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4626_ _0347_ _0369_ _0450_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_129_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4557_ _0345_ _0379_ _0380_ _0381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3508_ _1136_ _1675_ _1862_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_103_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4488_ _0310_ _0311_ _0312_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6227_ _2147_ _2186_ _2187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3439_ _1059_ _0839_ _1092_ _1103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_106_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6158_ _2065_ _2071_ _2110_ _2111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6227__A2 _2186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5109_ _0958_ _0959_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6089_ _2031_ _2035_ _2036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4410__A1 _0217_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4961__A2 _1949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5910__A1 _1537_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput30 net30 result[6] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_107_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6710__I0 _2663_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6716__S _2678_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5977__A1 _1612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6515__I _2264_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4401__A1 _0219_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3790_ _1598_ _2950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3874__I _3033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5460_ _1336_ _1343_ _1344_ _1346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4411_ _0231_ _0234_ _0235_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4704__A2 _0299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5901__A1 _1546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5391_ _1269_ _1270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4342_ _0102_ _2037_ _0166_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4273_ _0095_ _0096_ _0097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_114_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4468__A1 _3346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4468__B2 _3351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6012_ _3276_ _3278_ _1952_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
.ends

