magic
tech gf180mcuC
magscale 1 5
timestamp 1670060192
<< obsm1 >>
rect 672 1538 89320 58505
<< metal2 >>
rect 2464 59600 2520 60000
rect 6328 59600 6384 60000
rect 10192 59600 10248 60000
rect 14056 59600 14112 60000
rect 17920 59600 17976 60000
rect 21784 59600 21840 60000
rect 25648 59600 25704 60000
rect 29512 59600 29568 60000
rect 33376 59600 33432 60000
rect 37240 59600 37296 60000
rect 41104 59600 41160 60000
rect 44968 59600 45024 60000
rect 48832 59600 48888 60000
rect 52696 59600 52752 60000
rect 56560 59600 56616 60000
rect 60424 59600 60480 60000
rect 64288 59600 64344 60000
rect 68152 59600 68208 60000
rect 72016 59600 72072 60000
rect 75880 59600 75936 60000
rect 79744 59600 79800 60000
rect 83608 59600 83664 60000
rect 87472 59600 87528 60000
rect 4088 0 4144 400
rect 12264 0 12320 400
rect 20440 0 20496 400
rect 28616 0 28672 400
rect 36792 0 36848 400
rect 44968 0 45024 400
rect 53144 0 53200 400
rect 61320 0 61376 400
rect 69496 0 69552 400
rect 77672 0 77728 400
rect 85848 0 85904 400
<< obsm2 >>
rect 1806 59570 2434 59799
rect 2550 59570 6298 59799
rect 6414 59570 10162 59799
rect 10278 59570 14026 59799
rect 14142 59570 17890 59799
rect 18006 59570 21754 59799
rect 21870 59570 25618 59799
rect 25734 59570 29482 59799
rect 29598 59570 33346 59799
rect 33462 59570 37210 59799
rect 37326 59570 41074 59799
rect 41190 59570 44938 59799
rect 45054 59570 48802 59799
rect 48918 59570 52666 59799
rect 52782 59570 56530 59799
rect 56646 59570 60394 59799
rect 60510 59570 64258 59799
rect 64374 59570 68122 59799
rect 68238 59570 71986 59799
rect 72102 59570 75850 59799
rect 75966 59570 79714 59799
rect 79830 59570 83578 59799
rect 83694 59570 87442 59799
rect 87558 59570 87626 59799
rect 1806 430 87626 59570
rect 1806 400 4058 430
rect 4174 400 12234 430
rect 12350 400 20410 430
rect 20526 400 28586 430
rect 28702 400 36762 430
rect 36878 400 44938 430
rect 45054 400 53114 430
rect 53230 400 61290 430
rect 61406 400 69466 430
rect 69582 400 77642 430
rect 77758 400 85818 430
rect 85934 400 87626 430
<< obsm3 >>
rect 1801 1554 86855 59794
<< metal4 >>
rect 2224 1538 2384 58438
rect 9904 1538 10064 58438
rect 17584 1538 17744 58438
rect 25264 1538 25424 58438
rect 32944 1538 33104 58438
rect 40624 1538 40784 58438
rect 48304 1538 48464 58438
rect 55984 1538 56144 58438
rect 63664 1538 63824 58438
rect 71344 1538 71504 58438
rect 79024 1538 79184 58438
rect 86704 1538 86864 58438
<< obsm4 >>
rect 9422 58468 77882 59631
rect 9422 11489 9874 58468
rect 10094 11489 17554 58468
rect 17774 11489 25234 58468
rect 25454 11489 32914 58468
rect 33134 11489 40594 58468
rect 40814 11489 48274 58468
rect 48494 11489 55954 58468
rect 56174 11489 63634 58468
rect 63854 11489 71314 58468
rect 71534 11489 77882 58468
<< labels >>
rlabel metal2 s 75880 59600 75936 60000 6 Clock
port 1 nsew signal input
rlabel metal2 s 83608 59600 83664 60000 6 Enable
port 2 nsew signal input
rlabel metal2 s 4088 0 4144 400 6 K[0]
port 3 nsew signal input
rlabel metal2 s 12264 0 12320 400 6 K[1]
port 4 nsew signal input
rlabel metal2 s 20440 0 20496 400 6 K[2]
port 5 nsew signal input
rlabel metal2 s 2464 59600 2520 60000 6 Result[0]
port 6 nsew signal output
rlabel metal2 s 41104 59600 41160 60000 6 Result[10]
port 7 nsew signal output
rlabel metal2 s 44968 59600 45024 60000 6 Result[11]
port 8 nsew signal output
rlabel metal2 s 48832 59600 48888 60000 6 Result[12]
port 9 nsew signal output
rlabel metal2 s 52696 59600 52752 60000 6 Result[13]
port 10 nsew signal output
rlabel metal2 s 56560 59600 56616 60000 6 Result[14]
port 11 nsew signal output
rlabel metal2 s 60424 59600 60480 60000 6 Result[15]
port 12 nsew signal output
rlabel metal2 s 64288 59600 64344 60000 6 Result[16]
port 13 nsew signal output
rlabel metal2 s 6328 59600 6384 60000 6 Result[1]
port 14 nsew signal output
rlabel metal2 s 10192 59600 10248 60000 6 Result[2]
port 15 nsew signal output
rlabel metal2 s 14056 59600 14112 60000 6 Result[3]
port 16 nsew signal output
rlabel metal2 s 17920 59600 17976 60000 6 Result[4]
port 17 nsew signal output
rlabel metal2 s 21784 59600 21840 60000 6 Result[5]
port 18 nsew signal output
rlabel metal2 s 25648 59600 25704 60000 6 Result[6]
port 19 nsew signal output
rlabel metal2 s 29512 59600 29568 60000 6 Result[7]
port 20 nsew signal output
rlabel metal2 s 33376 59600 33432 60000 6 Result[8]
port 21 nsew signal output
rlabel metal2 s 37240 59600 37296 60000 6 Result[9]
port 22 nsew signal output
rlabel metal2 s 28616 0 28672 400 6 X[0]
port 23 nsew signal input
rlabel metal2 s 36792 0 36848 400 6 X[1]
port 24 nsew signal input
rlabel metal2 s 44968 0 45024 400 6 X[2]
port 25 nsew signal input
rlabel metal2 s 53144 0 53200 400 6 X[3]
port 26 nsew signal input
rlabel metal2 s 61320 0 61376 400 6 X[4]
port 27 nsew signal input
rlabel metal2 s 69496 0 69552 400 6 X[5]
port 28 nsew signal input
rlabel metal2 s 77672 0 77728 400 6 X[6]
port 29 nsew signal input
rlabel metal2 s 85848 0 85904 400 6 X[7]
port 30 nsew signal input
rlabel metal2 s 68152 59600 68208 60000 6 Z[0]
port 31 nsew signal input
rlabel metal2 s 72016 59600 72072 60000 6 Z[1]
port 32 nsew signal input
rlabel metal2 s 87472 59600 87528 60000 6 done
port 33 nsew signal output
rlabel metal2 s 79744 59600 79800 60000 6 reset
port 34 nsew signal input
rlabel metal4 s 2224 1538 2384 58438 6 vccd1
port 35 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 58438 6 vccd1
port 35 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 58438 6 vccd1
port 35 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 58438 6 vccd1
port 35 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 58438 6 vccd1
port 35 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 58438 6 vccd1
port 35 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 58438 6 vssd1
port 36 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 58438 6 vssd1
port 36 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 58438 6 vssd1
port 36 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 58438 6 vssd1
port 36 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 58438 6 vssd1
port 36 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 58438 6 vssd1
port 36 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 90000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 10863092
string GDS_FILE /home/radhe/tapeout_projects/radhe_gf180nm/openlane/multiply_komal/runs/22_12_03_15_03/results/signoff/multiply_komal.magic.gds
string GDS_START 449756
<< end >>

